
module pc_reg_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  XNOR2V2_8TH40 U1 ( .A1(A[31]), .A2(n28), .ZN(SUM[31]) );
  NAND2V2_8TH40 U2 ( .A1(n27), .A2(A[30]), .ZN(n28) );
  AND2V2_8TH40 U3 ( .A1(A[2]), .A2(A[3]), .Z(n1) );
  AND2V2_8TH40 U4 ( .A1(n1), .A2(A[4]), .Z(n2) );
  AND2V2_8TH40 U5 ( .A1(n2), .A2(A[5]), .Z(n3) );
  AND2V2_8TH40 U6 ( .A1(n3), .A2(A[6]), .Z(n4) );
  AND2V2_8TH40 U7 ( .A1(n4), .A2(A[7]), .Z(n5) );
  AND2V2_8TH40 U8 ( .A1(n5), .A2(A[8]), .Z(n6) );
  AND2V2_8TH40 U9 ( .A1(n6), .A2(A[9]), .Z(n7) );
  AND2V2_8TH40 U10 ( .A1(n7), .A2(A[10]), .Z(n8) );
  AND2V2_8TH40 U11 ( .A1(n8), .A2(A[11]), .Z(n9) );
  AND2V2_8TH40 U12 ( .A1(n9), .A2(A[12]), .Z(n10) );
  AND2V2_8TH40 U13 ( .A1(n10), .A2(A[13]), .Z(n11) );
  AND2V2_8TH40 U14 ( .A1(n11), .A2(A[14]), .Z(n12) );
  AND2V2_8TH40 U15 ( .A1(n12), .A2(A[15]), .Z(n13) );
  AND2V2_8TH40 U16 ( .A1(n13), .A2(A[16]), .Z(n14) );
  AND2V2_8TH40 U17 ( .A1(n14), .A2(A[17]), .Z(n15) );
  AND2V2_8TH40 U18 ( .A1(n15), .A2(A[18]), .Z(n16) );
  AND2V2_8TH40 U19 ( .A1(n16), .A2(A[19]), .Z(n17) );
  AND2V2_8TH40 U20 ( .A1(n17), .A2(A[20]), .Z(n18) );
  AND2V2_8TH40 U21 ( .A1(n18), .A2(A[21]), .Z(n19) );
  AND2V2_8TH40 U22 ( .A1(n19), .A2(A[22]), .Z(n20) );
  AND2V2_8TH40 U23 ( .A1(n20), .A2(A[23]), .Z(n21) );
  AND2V2_8TH40 U24 ( .A1(n21), .A2(A[24]), .Z(n22) );
  AND2V2_8TH40 U25 ( .A1(n22), .A2(A[25]), .Z(n23) );
  AND2V2_8TH40 U26 ( .A1(n23), .A2(A[26]), .Z(n24) );
  AND2V2_8TH40 U27 ( .A1(n24), .A2(A[27]), .Z(n25) );
  AND2V2_8TH40 U28 ( .A1(n25), .A2(A[28]), .Z(n26) );
  AND2V2_8TH40 U29 ( .A1(n26), .A2(A[29]), .Z(n27) );
  INV2_8TH40 U30 ( .I(A[2]), .ZN(SUM[2]) );
  XOR2V2_8TH40 U31 ( .A1(n27), .A2(A[30]), .Z(SUM[30]) );
  XOR2V2_8TH40 U32 ( .A1(n26), .A2(A[29]), .Z(SUM[29]) );
  XOR2V2_8TH40 U33 ( .A1(n25), .A2(A[28]), .Z(SUM[28]) );
  XOR2V2_8TH40 U34 ( .A1(n24), .A2(A[27]), .Z(SUM[27]) );
  XOR2V2_8TH40 U35 ( .A1(n23), .A2(A[26]), .Z(SUM[26]) );
  XOR2V2_8TH40 U36 ( .A1(n22), .A2(A[25]), .Z(SUM[25]) );
  XOR2V2_8TH40 U37 ( .A1(n21), .A2(A[24]), .Z(SUM[24]) );
  XOR2V2_8TH40 U38 ( .A1(n20), .A2(A[23]), .Z(SUM[23]) );
  XOR2V2_8TH40 U39 ( .A1(n19), .A2(A[22]), .Z(SUM[22]) );
  XOR2V2_8TH40 U40 ( .A1(n18), .A2(A[21]), .Z(SUM[21]) );
  XOR2V2_8TH40 U41 ( .A1(n17), .A2(A[20]), .Z(SUM[20]) );
  XOR2V2_8TH40 U42 ( .A1(n16), .A2(A[19]), .Z(SUM[19]) );
  XOR2V2_8TH40 U43 ( .A1(n15), .A2(A[18]), .Z(SUM[18]) );
  XOR2V2_8TH40 U44 ( .A1(n14), .A2(A[17]), .Z(SUM[17]) );
  XOR2V2_8TH40 U45 ( .A1(n13), .A2(A[16]), .Z(SUM[16]) );
  XOR2V2_8TH40 U46 ( .A1(n12), .A2(A[15]), .Z(SUM[15]) );
  XOR2V2_8TH40 U47 ( .A1(n11), .A2(A[14]), .Z(SUM[14]) );
  XOR2V2_8TH40 U48 ( .A1(n10), .A2(A[13]), .Z(SUM[13]) );
  XOR2V2_8TH40 U49 ( .A1(n9), .A2(A[12]), .Z(SUM[12]) );
  XOR2V2_8TH40 U50 ( .A1(n8), .A2(A[11]), .Z(SUM[11]) );
  XOR2V2_8TH40 U51 ( .A1(n7), .A2(A[10]), .Z(SUM[10]) );
  XOR2V2_8TH40 U52 ( .A1(n6), .A2(A[9]), .Z(SUM[9]) );
  XOR2V2_8TH40 U53 ( .A1(n5), .A2(A[8]), .Z(SUM[8]) );
  XOR2V2_8TH40 U54 ( .A1(n4), .A2(A[7]), .Z(SUM[7]) );
  XOR2V2_8TH40 U55 ( .A1(n3), .A2(A[6]), .Z(SUM[6]) );
  XOR2V2_8TH40 U56 ( .A1(n2), .A2(A[5]), .Z(SUM[5]) );
  XOR2V2_8TH40 U57 ( .A1(n1), .A2(A[4]), .Z(SUM[4]) );
  XOR2V2_8TH40 U58 ( .A1(A[2]), .A2(A[3]), .Z(SUM[3]) );
endmodule


module pc_reg ( clk, rst, stall_ctrl, branch_flag, branch_target_addr, pc_new, 
        pc, inst_mem_en, flush_BAR );
  input [5:0] stall_ctrl;
  input [31:0] branch_target_addr;
  input [31:0] pc_new;
  output [31:0] pc;
  input clk, rst, branch_flag, flush_BAR;
  output inst_mem_en;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21,
         N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71;

  DQV4_8TH40 inst_mem_en_reg ( .D(n71), .CK(clk), .Q(inst_mem_en) );
  DQV4_8TH40 pc_reg_0_ ( .D(n106), .CK(clk), .Q(pc[0]) );
  DQV4_8TH40 pc_reg_1_ ( .D(n105), .CK(clk), .Q(pc[1]) );
  DQV4_8TH40 pc_reg_2_ ( .D(n104), .CK(clk), .Q(pc[2]) );
  DQV4_8TH40 pc_reg_3_ ( .D(n103), .CK(clk), .Q(pc[3]) );
  DQV4_8TH40 pc_reg_4_ ( .D(n102), .CK(clk), .Q(pc[4]) );
  DQV4_8TH40 pc_reg_5_ ( .D(n101), .CK(clk), .Q(pc[5]) );
  DQV4_8TH40 pc_reg_6_ ( .D(n100), .CK(clk), .Q(pc[6]) );
  DQV4_8TH40 pc_reg_7_ ( .D(n99), .CK(clk), .Q(pc[7]) );
  DQV4_8TH40 pc_reg_8_ ( .D(n98), .CK(clk), .Q(pc[8]) );
  DQV4_8TH40 pc_reg_9_ ( .D(n97), .CK(clk), .Q(pc[9]) );
  DQV4_8TH40 pc_reg_10_ ( .D(n96), .CK(clk), .Q(pc[10]) );
  DQV4_8TH40 pc_reg_11_ ( .D(n95), .CK(clk), .Q(pc[11]) );
  DQV4_8TH40 pc_reg_12_ ( .D(n94), .CK(clk), .Q(pc[12]) );
  DQV4_8TH40 pc_reg_13_ ( .D(n93), .CK(clk), .Q(pc[13]) );
  DQV4_8TH40 pc_reg_14_ ( .D(n92), .CK(clk), .Q(pc[14]) );
  DQV4_8TH40 pc_reg_15_ ( .D(n91), .CK(clk), .Q(pc[15]) );
  DQV4_8TH40 pc_reg_16_ ( .D(n90), .CK(clk), .Q(pc[16]) );
  DQV4_8TH40 pc_reg_17_ ( .D(n89), .CK(clk), .Q(pc[17]) );
  DQV4_8TH40 pc_reg_18_ ( .D(n88), .CK(clk), .Q(pc[18]) );
  DQV4_8TH40 pc_reg_19_ ( .D(n87), .CK(clk), .Q(pc[19]) );
  DQV4_8TH40 pc_reg_20_ ( .D(n86), .CK(clk), .Q(pc[20]) );
  DQV4_8TH40 pc_reg_21_ ( .D(n85), .CK(clk), .Q(pc[21]) );
  DQV4_8TH40 pc_reg_22_ ( .D(n84), .CK(clk), .Q(pc[22]) );
  DQV4_8TH40 pc_reg_23_ ( .D(n83), .CK(clk), .Q(pc[23]) );
  DQV4_8TH40 pc_reg_24_ ( .D(n82), .CK(clk), .Q(pc[24]) );
  DQV4_8TH40 pc_reg_25_ ( .D(n81), .CK(clk), .Q(pc[25]) );
  DQV4_8TH40 pc_reg_26_ ( .D(n80), .CK(clk), .Q(pc[26]) );
  DQV4_8TH40 pc_reg_27_ ( .D(n79), .CK(clk), .Q(pc[27]) );
  DQV4_8TH40 pc_reg_28_ ( .D(n78), .CK(clk), .Q(pc[28]) );
  DQV4_8TH40 pc_reg_29_ ( .D(n77), .CK(clk), .Q(pc[29]) );
  DQV4_8TH40 pc_reg_30_ ( .D(n76), .CK(clk), .Q(pc[30]) );
  DQV4_8TH40 pc_reg_31_ ( .D(n75), .CK(clk), .Q(pc[31]) );
  pc_reg_DW01_add_0 add_41 ( .A(pc), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, N10, N9, N8}) );
  NAND2V2_8TH40 U3 ( .A1(n54), .A2(n55), .ZN(n75) );
  AOI22V2_8TH40 U4 ( .A1(branch_target_addr[31]), .A2(n6), .B1(pc[31]), .B2(n7), .ZN(n54) );
  NAND2V2_8TH40 U6 ( .A1(n52), .A2(n53), .ZN(n76) );
  AOI22V2_8TH40 U7 ( .A1(branch_target_addr[30]), .A2(n6), .B1(pc[30]), .B2(n7), .ZN(n52) );
  NAND2V2_8TH40 U8 ( .A1(n50), .A2(n51), .ZN(n77) );
  AOI22V2_8TH40 U9 ( .A1(branch_target_addr[29]), .A2(n6), .B1(pc[29]), .B2(n7), .ZN(n50) );
  NAND2V2_8TH40 U10 ( .A1(n48), .A2(n49), .ZN(n78) );
  AOI22V2_8TH40 U11 ( .A1(branch_target_addr[28]), .A2(n6), .B1(pc[28]), .B2(
        n7), .ZN(n48) );
  NAND2V2_8TH40 U12 ( .A1(n46), .A2(n47), .ZN(n79) );
  AOI22V2_8TH40 U13 ( .A1(branch_target_addr[27]), .A2(n6), .B1(pc[27]), .B2(
        n7), .ZN(n46) );
  NAND2V2_8TH40 U14 ( .A1(n44), .A2(n45), .ZN(n80) );
  AOI22V2_8TH40 U15 ( .A1(branch_target_addr[26]), .A2(n6), .B1(pc[26]), .B2(
        n7), .ZN(n44) );
  NAND2V2_8TH40 U16 ( .A1(n42), .A2(n43), .ZN(n81) );
  AOI22V2_8TH40 U17 ( .A1(branch_target_addr[25]), .A2(n6), .B1(pc[25]), .B2(
        n7), .ZN(n42) );
  NAND2V2_8TH40 U18 ( .A1(n40), .A2(n41), .ZN(n82) );
  AOI22V2_8TH40 U19 ( .A1(branch_target_addr[24]), .A2(n6), .B1(pc[24]), .B2(
        n7), .ZN(n40) );
  NAND2V2_8TH40 U20 ( .A1(n38), .A2(n39), .ZN(n83) );
  AOI22V2_8TH40 U21 ( .A1(branch_target_addr[23]), .A2(n6), .B1(pc[23]), .B2(
        n7), .ZN(n38) );
  NAND2V2_8TH40 U22 ( .A1(n36), .A2(n37), .ZN(n84) );
  AOI22V2_8TH40 U23 ( .A1(branch_target_addr[22]), .A2(n6), .B1(pc[22]), .B2(
        n7), .ZN(n36) );
  NAND2V2_8TH40 U24 ( .A1(n34), .A2(n35), .ZN(n85) );
  AOI22V2_8TH40 U25 ( .A1(branch_target_addr[21]), .A2(n6), .B1(pc[21]), .B2(
        n7), .ZN(n34) );
  NAND2V2_8TH40 U26 ( .A1(n32), .A2(n33), .ZN(n86) );
  AOI22V2_8TH40 U27 ( .A1(branch_target_addr[20]), .A2(n6), .B1(pc[20]), .B2(
        n7), .ZN(n32) );
  NAND2V2_8TH40 U28 ( .A1(n30), .A2(n31), .ZN(n87) );
  AOI22V2_8TH40 U29 ( .A1(branch_target_addr[19]), .A2(n6), .B1(pc[19]), .B2(
        n7), .ZN(n30) );
  NAND2V2_8TH40 U30 ( .A1(n28), .A2(n29), .ZN(n88) );
  AOI22V2_8TH40 U31 ( .A1(branch_target_addr[18]), .A2(n6), .B1(pc[18]), .B2(
        n7), .ZN(n28) );
  NAND2V2_8TH40 U32 ( .A1(n26), .A2(n27), .ZN(n89) );
  AOI22V2_8TH40 U33 ( .A1(branch_target_addr[17]), .A2(n6), .B1(pc[17]), .B2(
        n7), .ZN(n26) );
  NAND2V2_8TH40 U34 ( .A1(n24), .A2(n25), .ZN(n90) );
  AOI22V2_8TH40 U35 ( .A1(branch_target_addr[16]), .A2(n6), .B1(pc[16]), .B2(
        n7), .ZN(n24) );
  NAND2V2_8TH40 U36 ( .A1(n22), .A2(n23), .ZN(n91) );
  AOI22V2_8TH40 U37 ( .A1(branch_target_addr[15]), .A2(n6), .B1(pc[15]), .B2(
        n7), .ZN(n22) );
  NAND2V2_8TH40 U38 ( .A1(n20), .A2(n21), .ZN(n92) );
  AOI22V2_8TH40 U39 ( .A1(branch_target_addr[14]), .A2(n6), .B1(pc[14]), .B2(
        n7), .ZN(n20) );
  NAND2V2_8TH40 U40 ( .A1(n18), .A2(n19), .ZN(n93) );
  AOI22V2_8TH40 U41 ( .A1(branch_target_addr[13]), .A2(n6), .B1(pc[13]), .B2(
        n7), .ZN(n18) );
  NAND2V2_8TH40 U42 ( .A1(n16), .A2(n17), .ZN(n94) );
  AOI22V2_8TH40 U43 ( .A1(branch_target_addr[12]), .A2(n6), .B1(pc[12]), .B2(
        n7), .ZN(n16) );
  NAND2V2_8TH40 U44 ( .A1(n14), .A2(n15), .ZN(n95) );
  AOI22V2_8TH40 U45 ( .A1(branch_target_addr[11]), .A2(n6), .B1(pc[11]), .B2(
        n7), .ZN(n14) );
  NAND2V2_8TH40 U46 ( .A1(n12), .A2(n13), .ZN(n96) );
  AOI22V2_8TH40 U47 ( .A1(branch_target_addr[10]), .A2(n6), .B1(pc[10]), .B2(
        n7), .ZN(n12) );
  NAND2V2_8TH40 U48 ( .A1(n10), .A2(n11), .ZN(n97) );
  AOI22V2_8TH40 U49 ( .A1(branch_target_addr[9]), .A2(n6), .B1(pc[9]), .B2(n7), 
        .ZN(n10) );
  NAND2V2_8TH40 U50 ( .A1(n8), .A2(n9), .ZN(n98) );
  AOI22V2_8TH40 U51 ( .A1(branch_target_addr[8]), .A2(n6), .B1(pc[8]), .B2(n7), 
        .ZN(n8) );
  NAND2V2_8TH40 U52 ( .A1(n2), .A2(n3), .ZN(n99) );
  AOI22V2_8TH40 U53 ( .A1(branch_target_addr[7]), .A2(n6), .B1(pc[7]), .B2(n7), 
        .ZN(n2) );
  NAND2V2_8TH40 U54 ( .A1(n68), .A2(n69), .ZN(n100) );
  AOI22V2_8TH40 U55 ( .A1(branch_target_addr[6]), .A2(n6), .B1(pc[6]), .B2(n7), 
        .ZN(n68) );
  NAND2V2_8TH40 U56 ( .A1(n66), .A2(n67), .ZN(n101) );
  AOI22V2_8TH40 U57 ( .A1(branch_target_addr[5]), .A2(n6), .B1(pc[5]), .B2(n7), 
        .ZN(n66) );
  NAND2V2_8TH40 U58 ( .A1(n64), .A2(n65), .ZN(n102) );
  AOI22V2_8TH40 U59 ( .A1(branch_target_addr[4]), .A2(n6), .B1(pc[4]), .B2(n7), 
        .ZN(n64) );
  NAND2V2_8TH40 U60 ( .A1(n62), .A2(n63), .ZN(n103) );
  AOI22V2_8TH40 U61 ( .A1(branch_target_addr[3]), .A2(n6), .B1(pc[3]), .B2(n7), 
        .ZN(n62) );
  AOI22V2_8TH40 U62 ( .A1(N11), .A2(n4), .B1(pc_new[3]), .B2(n5), .ZN(n63) );
  NAND2V2_8TH40 U63 ( .A1(n60), .A2(n61), .ZN(n104) );
  AOI22V2_8TH40 U64 ( .A1(branch_target_addr[2]), .A2(n6), .B1(pc[2]), .B2(n7), 
        .ZN(n60) );
  AOI22V2_8TH40 U65 ( .A1(N10), .A2(n4), .B1(pc_new[2]), .B2(n5), .ZN(n61) );
  NAND2V2_8TH40 U66 ( .A1(n58), .A2(n59), .ZN(n105) );
  AOI22V2_8TH40 U67 ( .A1(branch_target_addr[1]), .A2(n6), .B1(pc[1]), .B2(n7), 
        .ZN(n58) );
  AOI22V2_8TH40 U68 ( .A1(N9), .A2(n4), .B1(pc_new[1]), .B2(n5), .ZN(n59) );
  NAND2V2_8TH40 U69 ( .A1(n56), .A2(n57), .ZN(n106) );
  AOI22V2_8TH40 U70 ( .A1(branch_target_addr[0]), .A2(n6), .B1(pc[0]), .B2(n7), 
        .ZN(n56) );
  AOI22V2_8TH40 U71 ( .A1(N8), .A2(n4), .B1(pc_new[0]), .B2(n5), .ZN(n57) );
  CLKNV1_8TH40 U72 ( .I(rst), .ZN(n71) );
  AOI22V0_8TH40 U73 ( .A1(N15), .A2(n4), .B1(pc_new[7]), .B2(n5), .ZN(n3) );
  AOI22V0_8TH40 U74 ( .A1(N16), .A2(n4), .B1(pc_new[8]), .B2(n5), .ZN(n9) );
  AOI22V0_8TH40 U75 ( .A1(N17), .A2(n4), .B1(pc_new[9]), .B2(n5), .ZN(n11) );
  AOI22V0_8TH40 U76 ( .A1(N18), .A2(n4), .B1(pc_new[10]), .B2(n5), .ZN(n13) );
  AOI22V0_8TH40 U77 ( .A1(N19), .A2(n4), .B1(pc_new[11]), .B2(n5), .ZN(n15) );
  AOI22V0_8TH40 U78 ( .A1(N20), .A2(n4), .B1(pc_new[12]), .B2(n5), .ZN(n17) );
  AOI22V0_8TH40 U79 ( .A1(N21), .A2(n4), .B1(pc_new[13]), .B2(n5), .ZN(n19) );
  AOI22V0_8TH40 U80 ( .A1(N22), .A2(n4), .B1(pc_new[14]), .B2(n5), .ZN(n21) );
  AOI22V0_8TH40 U81 ( .A1(N23), .A2(n4), .B1(pc_new[15]), .B2(n5), .ZN(n23) );
  AOI22V0_8TH40 U82 ( .A1(N24), .A2(n4), .B1(pc_new[16]), .B2(n5), .ZN(n25) );
  AOI22V0_8TH40 U83 ( .A1(N25), .A2(n4), .B1(pc_new[17]), .B2(n5), .ZN(n27) );
  AOI22V0_8TH40 U84 ( .A1(N26), .A2(n4), .B1(pc_new[18]), .B2(n5), .ZN(n29) );
  AOI22V0_8TH40 U85 ( .A1(N27), .A2(n4), .B1(pc_new[19]), .B2(n5), .ZN(n31) );
  AOI22V0_8TH40 U86 ( .A1(N28), .A2(n4), .B1(pc_new[20]), .B2(n5), .ZN(n33) );
  AOI22V0_8TH40 U87 ( .A1(N29), .A2(n4), .B1(pc_new[21]), .B2(n5), .ZN(n35) );
  AOI22V0_8TH40 U88 ( .A1(N30), .A2(n4), .B1(pc_new[22]), .B2(n5), .ZN(n37) );
  AOI22V0_8TH40 U89 ( .A1(N31), .A2(n4), .B1(pc_new[23]), .B2(n5), .ZN(n39) );
  AOI22V0_8TH40 U90 ( .A1(N32), .A2(n4), .B1(pc_new[24]), .B2(n5), .ZN(n41) );
  AOI22V0_8TH40 U91 ( .A1(N33), .A2(n4), .B1(pc_new[25]), .B2(n5), .ZN(n43) );
  AOI22V0_8TH40 U92 ( .A1(N34), .A2(n4), .B1(pc_new[26]), .B2(n5), .ZN(n45) );
  AOI22V0_8TH40 U93 ( .A1(N35), .A2(n4), .B1(pc_new[27]), .B2(n5), .ZN(n47) );
  AOI22V0_8TH40 U94 ( .A1(N36), .A2(n4), .B1(pc_new[28]), .B2(n5), .ZN(n49) );
  AOI22V0_8TH40 U95 ( .A1(N37), .A2(n4), .B1(pc_new[29]), .B2(n5), .ZN(n51) );
  AOI22V0_8TH40 U96 ( .A1(N38), .A2(n4), .B1(pc_new[30]), .B2(n5), .ZN(n53) );
  AOI22V0_8TH40 U97 ( .A1(N39), .A2(n4), .B1(pc_new[31]), .B2(n5), .ZN(n55) );
  AOI22V0_8TH40 U98 ( .A1(N12), .A2(n4), .B1(pc_new[4]), .B2(n5), .ZN(n65) );
  AOI22V0_8TH40 U99 ( .A1(N13), .A2(n4), .B1(pc_new[5]), .B2(n5), .ZN(n67) );
  AOI22V0_8TH40 U100 ( .A1(N14), .A2(n4), .B1(pc_new[6]), .B2(n5), .ZN(n69) );
  INOR2V0_8TH40 U101 ( .A1(inst_mem_en), .B1(flush_BAR), .ZN(n5) );
  I2NOR4V0_8TH40 U102 ( .A1(inst_mem_en), .A2(flush_BAR), .B1(n7), .B2(
        branch_flag), .ZN(n4) );
  CLKNV1_8TH40 U103 ( .I(n70), .ZN(n7) );
  AND4V0_8TH40 U104 ( .A1(branch_flag), .A2(inst_mem_en), .A3(flush_BAR), .A4(
        n70), .Z(n6) );
  NAND3V0P5_8TH40 U105 ( .A1(inst_mem_en), .A2(flush_BAR), .A3(stall_ctrl[0]), 
        .ZN(n70) );
endmodule


module pipe_reg_ifid ( clk, rst, stall_ctrl, if_pc, if_inst, id_pc, id_inst, 
        flush_BAR );
  input [5:0] stall_ctrl;
  input [31:0] if_pc;
  input [31:0] if_inst;
  output [31:0] id_pc;
  output [31:0] id_inst;
  input clk, rst, flush_BAR;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n1, n2, n3, n68;

  DQV4_8TH40 id_inst_reg_31_ ( .D(n67), .CK(clk), .Q(id_inst[31]) );
  DQV4_8TH40 id_inst_reg_30_ ( .D(n66), .CK(clk), .Q(id_inst[30]) );
  DQV4_8TH40 id_inst_reg_29_ ( .D(n65), .CK(clk), .Q(id_inst[29]) );
  DQV4_8TH40 id_inst_reg_28_ ( .D(n64), .CK(clk), .Q(id_inst[28]) );
  DQV4_8TH40 id_inst_reg_27_ ( .D(n63), .CK(clk), .Q(id_inst[27]) );
  DQV4_8TH40 id_inst_reg_26_ ( .D(n62), .CK(clk), .Q(id_inst[26]) );
  DQV4_8TH40 id_inst_reg_25_ ( .D(n61), .CK(clk), .Q(id_inst[25]) );
  DQV4_8TH40 id_inst_reg_24_ ( .D(n60), .CK(clk), .Q(id_inst[24]) );
  DQV4_8TH40 id_inst_reg_23_ ( .D(n59), .CK(clk), .Q(id_inst[23]) );
  DQV4_8TH40 id_inst_reg_22_ ( .D(n58), .CK(clk), .Q(id_inst[22]) );
  DQV4_8TH40 id_inst_reg_21_ ( .D(n57), .CK(clk), .Q(id_inst[21]) );
  DQV4_8TH40 id_inst_reg_20_ ( .D(n56), .CK(clk), .Q(id_inst[20]) );
  DQV4_8TH40 id_inst_reg_19_ ( .D(n55), .CK(clk), .Q(id_inst[19]) );
  DQV4_8TH40 id_inst_reg_18_ ( .D(n54), .CK(clk), .Q(id_inst[18]) );
  DQV4_8TH40 id_inst_reg_17_ ( .D(n53), .CK(clk), .Q(id_inst[17]) );
  DQV4_8TH40 id_inst_reg_16_ ( .D(n52), .CK(clk), .Q(id_inst[16]) );
  DQV4_8TH40 id_inst_reg_15_ ( .D(n51), .CK(clk), .Q(id_inst[15]) );
  DQV4_8TH40 id_inst_reg_14_ ( .D(n50), .CK(clk), .Q(id_inst[14]) );
  DQV4_8TH40 id_inst_reg_13_ ( .D(n49), .CK(clk), .Q(id_inst[13]) );
  DQV4_8TH40 id_inst_reg_12_ ( .D(n48), .CK(clk), .Q(id_inst[12]) );
  DQV4_8TH40 id_inst_reg_11_ ( .D(n47), .CK(clk), .Q(id_inst[11]) );
  DQV4_8TH40 id_inst_reg_10_ ( .D(n46), .CK(clk), .Q(id_inst[10]) );
  DQV4_8TH40 id_inst_reg_9_ ( .D(n45), .CK(clk), .Q(id_inst[9]) );
  DQV4_8TH40 id_inst_reg_8_ ( .D(n44), .CK(clk), .Q(id_inst[8]) );
  DQV4_8TH40 id_inst_reg_7_ ( .D(n43), .CK(clk), .Q(id_inst[7]) );
  DQV4_8TH40 id_inst_reg_6_ ( .D(n42), .CK(clk), .Q(id_inst[6]) );
  DQV4_8TH40 id_inst_reg_5_ ( .D(n41), .CK(clk), .Q(id_inst[5]) );
  DQV4_8TH40 id_inst_reg_4_ ( .D(n40), .CK(clk), .Q(id_inst[4]) );
  DQV4_8TH40 id_inst_reg_3_ ( .D(n39), .CK(clk), .Q(id_inst[3]) );
  DQV4_8TH40 id_inst_reg_2_ ( .D(n38), .CK(clk), .Q(id_inst[2]) );
  DQV4_8TH40 id_inst_reg_1_ ( .D(n37), .CK(clk), .Q(id_inst[1]) );
  DQV4_8TH40 id_inst_reg_0_ ( .D(n36), .CK(clk), .Q(id_inst[0]) );
  DQV4_8TH40 id_pc_reg_31_ ( .D(n35), .CK(clk), .Q(id_pc[31]) );
  DQV4_8TH40 id_pc_reg_30_ ( .D(n34), .CK(clk), .Q(id_pc[30]) );
  DQV4_8TH40 id_pc_reg_29_ ( .D(n33), .CK(clk), .Q(id_pc[29]) );
  DQV4_8TH40 id_pc_reg_28_ ( .D(n32), .CK(clk), .Q(id_pc[28]) );
  DQV4_8TH40 id_pc_reg_27_ ( .D(n31), .CK(clk), .Q(id_pc[27]) );
  DQV4_8TH40 id_pc_reg_26_ ( .D(n30), .CK(clk), .Q(id_pc[26]) );
  DQV4_8TH40 id_pc_reg_25_ ( .D(n29), .CK(clk), .Q(id_pc[25]) );
  DQV4_8TH40 id_pc_reg_24_ ( .D(n28), .CK(clk), .Q(id_pc[24]) );
  DQV4_8TH40 id_pc_reg_23_ ( .D(n27), .CK(clk), .Q(id_pc[23]) );
  DQV4_8TH40 id_pc_reg_22_ ( .D(n26), .CK(clk), .Q(id_pc[22]) );
  DQV4_8TH40 id_pc_reg_21_ ( .D(n25), .CK(clk), .Q(id_pc[21]) );
  DQV4_8TH40 id_pc_reg_20_ ( .D(n24), .CK(clk), .Q(id_pc[20]) );
  DQV4_8TH40 id_pc_reg_19_ ( .D(n23), .CK(clk), .Q(id_pc[19]) );
  DQV4_8TH40 id_pc_reg_18_ ( .D(n22), .CK(clk), .Q(id_pc[18]) );
  DQV4_8TH40 id_pc_reg_17_ ( .D(n21), .CK(clk), .Q(id_pc[17]) );
  DQV4_8TH40 id_pc_reg_16_ ( .D(n20), .CK(clk), .Q(id_pc[16]) );
  DQV4_8TH40 id_pc_reg_15_ ( .D(n19), .CK(clk), .Q(id_pc[15]) );
  DQV4_8TH40 id_pc_reg_14_ ( .D(n18), .CK(clk), .Q(id_pc[14]) );
  DQV4_8TH40 id_pc_reg_13_ ( .D(n17), .CK(clk), .Q(id_pc[13]) );
  DQV4_8TH40 id_pc_reg_12_ ( .D(n16), .CK(clk), .Q(id_pc[12]) );
  DQV4_8TH40 id_pc_reg_11_ ( .D(n15), .CK(clk), .Q(id_pc[11]) );
  DQV4_8TH40 id_pc_reg_10_ ( .D(n14), .CK(clk), .Q(id_pc[10]) );
  DQV4_8TH40 id_pc_reg_9_ ( .D(n13), .CK(clk), .Q(id_pc[9]) );
  DQV4_8TH40 id_pc_reg_8_ ( .D(n12), .CK(clk), .Q(id_pc[8]) );
  DQV4_8TH40 id_pc_reg_7_ ( .D(n11), .CK(clk), .Q(id_pc[7]) );
  DQV4_8TH40 id_pc_reg_6_ ( .D(n10), .CK(clk), .Q(id_pc[6]) );
  DQV4_8TH40 id_pc_reg_5_ ( .D(n9), .CK(clk), .Q(id_pc[5]) );
  DQV4_8TH40 id_pc_reg_4_ ( .D(n8), .CK(clk), .Q(id_pc[4]) );
  DQV4_8TH40 id_pc_reg_3_ ( .D(n7), .CK(clk), .Q(id_pc[3]) );
  DQV4_8TH40 id_pc_reg_2_ ( .D(n6), .CK(clk), .Q(id_pc[2]) );
  DQV4_8TH40 id_pc_reg_1_ ( .D(n5), .CK(clk), .Q(id_pc[1]) );
  DQV4_8TH40 id_pc_reg_0_ ( .D(n4), .CK(clk), .Q(id_pc[0]) );
  INV2_8TH40 U2 ( .I(n68), .ZN(n1) );
  INV2_8TH40 U3 ( .I(n1), .ZN(n2) );
  INOR3V0_8TH40 U4 ( .A1(flush_BAR), .B1(n3), .B2(rst), .ZN(n68) );
  AO22V4_8TH40 U5 ( .A1(id_inst[31]), .A2(n3), .B1(if_inst[31]), .B2(n2), .Z(
        n67) );
  AO22V4_8TH40 U6 ( .A1(id_inst[30]), .A2(n3), .B1(if_inst[30]), .B2(n2), .Z(
        n66) );
  AO22V4_8TH40 U7 ( .A1(id_inst[29]), .A2(n3), .B1(if_inst[29]), .B2(n2), .Z(
        n65) );
  AO22V4_8TH40 U8 ( .A1(id_inst[28]), .A2(n3), .B1(if_inst[28]), .B2(n2), .Z(
        n64) );
  AO22V4_8TH40 U9 ( .A1(id_inst[27]), .A2(n3), .B1(if_inst[27]), .B2(n2), .Z(
        n63) );
  AO22V4_8TH40 U10 ( .A1(id_inst[26]), .A2(n3), .B1(if_inst[26]), .B2(n2), .Z(
        n62) );
  AO22V4_8TH40 U11 ( .A1(id_inst[25]), .A2(n3), .B1(if_inst[25]), .B2(n2), .Z(
        n61) );
  AO22V4_8TH40 U12 ( .A1(id_inst[24]), .A2(n3), .B1(if_inst[24]), .B2(n2), .Z(
        n60) );
  AO22V4_8TH40 U13 ( .A1(id_inst[23]), .A2(n3), .B1(if_inst[23]), .B2(n2), .Z(
        n59) );
  AO22V4_8TH40 U14 ( .A1(id_inst[22]), .A2(n3), .B1(if_inst[22]), .B2(n2), .Z(
        n58) );
  AO22V4_8TH40 U15 ( .A1(id_inst[21]), .A2(n3), .B1(if_inst[21]), .B2(n2), .Z(
        n57) );
  AO22V4_8TH40 U16 ( .A1(id_inst[20]), .A2(n3), .B1(if_inst[20]), .B2(n2), .Z(
        n56) );
  AO22V4_8TH40 U17 ( .A1(id_inst[19]), .A2(n3), .B1(if_inst[19]), .B2(n2), .Z(
        n55) );
  AO22V4_8TH40 U18 ( .A1(id_inst[18]), .A2(n3), .B1(if_inst[18]), .B2(n2), .Z(
        n54) );
  AO22V4_8TH40 U19 ( .A1(id_inst[17]), .A2(n3), .B1(if_inst[17]), .B2(n2), .Z(
        n53) );
  AO22V4_8TH40 U20 ( .A1(id_inst[16]), .A2(n3), .B1(if_inst[16]), .B2(n2), .Z(
        n52) );
  AO22V4_8TH40 U21 ( .A1(id_inst[15]), .A2(n3), .B1(if_inst[15]), .B2(n2), .Z(
        n51) );
  AO22V4_8TH40 U22 ( .A1(id_inst[14]), .A2(n3), .B1(if_inst[14]), .B2(n2), .Z(
        n50) );
  AO22V4_8TH40 U23 ( .A1(id_inst[13]), .A2(n3), .B1(if_inst[13]), .B2(n2), .Z(
        n49) );
  AO22V4_8TH40 U24 ( .A1(id_inst[12]), .A2(n3), .B1(if_inst[12]), .B2(n2), .Z(
        n48) );
  AO22V4_8TH40 U25 ( .A1(id_inst[11]), .A2(n3), .B1(if_inst[11]), .B2(n2), .Z(
        n47) );
  AO22V4_8TH40 U26 ( .A1(id_inst[10]), .A2(n3), .B1(if_inst[10]), .B2(n2), .Z(
        n46) );
  AO22V4_8TH40 U27 ( .A1(id_inst[9]), .A2(n3), .B1(if_inst[9]), .B2(n2), .Z(
        n45) );
  AO22V4_8TH40 U28 ( .A1(id_inst[8]), .A2(n3), .B1(if_inst[8]), .B2(n2), .Z(
        n44) );
  AO22V4_8TH40 U29 ( .A1(id_inst[7]), .A2(n3), .B1(if_inst[7]), .B2(n2), .Z(
        n43) );
  AO22V4_8TH40 U30 ( .A1(id_inst[6]), .A2(n3), .B1(if_inst[6]), .B2(n2), .Z(
        n42) );
  AO22V4_8TH40 U31 ( .A1(id_inst[5]), .A2(n3), .B1(if_inst[5]), .B2(n2), .Z(
        n41) );
  AO22V4_8TH40 U32 ( .A1(id_inst[4]), .A2(n3), .B1(if_inst[4]), .B2(n2), .Z(
        n40) );
  AO22V4_8TH40 U33 ( .A1(id_inst[3]), .A2(n3), .B1(if_inst[3]), .B2(n2), .Z(
        n39) );
  AO22V4_8TH40 U34 ( .A1(id_inst[2]), .A2(n3), .B1(if_inst[2]), .B2(n2), .Z(
        n38) );
  AO22V4_8TH40 U35 ( .A1(id_inst[1]), .A2(n3), .B1(if_inst[1]), .B2(n2), .Z(
        n37) );
  AO22V4_8TH40 U36 ( .A1(id_inst[0]), .A2(n3), .B1(if_inst[0]), .B2(n2), .Z(
        n36) );
  AO22V0_8TH40 U37 ( .A1(id_pc[5]), .A2(n3), .B1(if_pc[5]), .B2(n2), .Z(n9) );
  AO22V0_8TH40 U38 ( .A1(id_pc[4]), .A2(n3), .B1(if_pc[4]), .B2(n2), .Z(n8) );
  AO22V0_8TH40 U39 ( .A1(id_pc[3]), .A2(n3), .B1(if_pc[3]), .B2(n2), .Z(n7) );
  AO22V0_8TH40 U40 ( .A1(id_pc[2]), .A2(n3), .B1(if_pc[2]), .B2(n2), .Z(n6) );
  AO22V0_8TH40 U41 ( .A1(id_pc[1]), .A2(n3), .B1(if_pc[1]), .B2(n2), .Z(n5) );
  AO22V0_8TH40 U42 ( .A1(id_pc[0]), .A2(n3), .B1(if_pc[0]), .B2(n2), .Z(n4) );
  AO22V0_8TH40 U43 ( .A1(id_pc[31]), .A2(n3), .B1(if_pc[31]), .B2(n2), .Z(n35)
         );
  AO22V0_8TH40 U44 ( .A1(id_pc[30]), .A2(n3), .B1(if_pc[30]), .B2(n2), .Z(n34)
         );
  AO22V0_8TH40 U45 ( .A1(id_pc[29]), .A2(n3), .B1(if_pc[29]), .B2(n2), .Z(n33)
         );
  AO22V0_8TH40 U46 ( .A1(id_pc[28]), .A2(n3), .B1(if_pc[28]), .B2(n2), .Z(n32)
         );
  AO22V0_8TH40 U47 ( .A1(id_pc[27]), .A2(n3), .B1(if_pc[27]), .B2(n2), .Z(n31)
         );
  AO22V0_8TH40 U48 ( .A1(id_pc[26]), .A2(n3), .B1(if_pc[26]), .B2(n2), .Z(n30)
         );
  AO22V0_8TH40 U49 ( .A1(id_pc[25]), .A2(n3), .B1(if_pc[25]), .B2(n2), .Z(n29)
         );
  AO22V0_8TH40 U50 ( .A1(id_pc[24]), .A2(n3), .B1(if_pc[24]), .B2(n2), .Z(n28)
         );
  AO22V0_8TH40 U51 ( .A1(id_pc[23]), .A2(n3), .B1(if_pc[23]), .B2(n2), .Z(n27)
         );
  AO22V0_8TH40 U52 ( .A1(id_pc[22]), .A2(n3), .B1(if_pc[22]), .B2(n2), .Z(n26)
         );
  AO22V0_8TH40 U53 ( .A1(id_pc[21]), .A2(n3), .B1(if_pc[21]), .B2(n2), .Z(n25)
         );
  AO22V0_8TH40 U54 ( .A1(id_pc[20]), .A2(n3), .B1(if_pc[20]), .B2(n2), .Z(n24)
         );
  AO22V0_8TH40 U55 ( .A1(id_pc[19]), .A2(n3), .B1(if_pc[19]), .B2(n2), .Z(n23)
         );
  AO22V0_8TH40 U56 ( .A1(id_pc[18]), .A2(n3), .B1(if_pc[18]), .B2(n2), .Z(n22)
         );
  AO22V0_8TH40 U57 ( .A1(id_pc[17]), .A2(n3), .B1(if_pc[17]), .B2(n2), .Z(n21)
         );
  AO22V0_8TH40 U58 ( .A1(id_pc[16]), .A2(n3), .B1(if_pc[16]), .B2(n2), .Z(n20)
         );
  AO22V0_8TH40 U59 ( .A1(id_pc[15]), .A2(n3), .B1(if_pc[15]), .B2(n2), .Z(n19)
         );
  AO22V0_8TH40 U60 ( .A1(id_pc[14]), .A2(n3), .B1(if_pc[14]), .B2(n2), .Z(n18)
         );
  AO22V0_8TH40 U61 ( .A1(id_pc[13]), .A2(n3), .B1(if_pc[13]), .B2(n2), .Z(n17)
         );
  AO22V0_8TH40 U62 ( .A1(id_pc[12]), .A2(n3), .B1(if_pc[12]), .B2(n2), .Z(n16)
         );
  AO22V0_8TH40 U63 ( .A1(id_pc[11]), .A2(n3), .B1(if_pc[11]), .B2(n2), .Z(n15)
         );
  AO22V0_8TH40 U64 ( .A1(id_pc[10]), .A2(n3), .B1(if_pc[10]), .B2(n2), .Z(n14)
         );
  AO22V0_8TH40 U65 ( .A1(id_pc[9]), .A2(n3), .B1(if_pc[9]), .B2(n2), .Z(n13)
         );
  AO22V0_8TH40 U66 ( .A1(id_pc[8]), .A2(n3), .B1(if_pc[8]), .B2(n2), .Z(n12)
         );
  AO22V0_8TH40 U67 ( .A1(id_pc[7]), .A2(n3), .B1(if_pc[7]), .B2(n2), .Z(n11)
         );
  AO22V0_8TH40 U68 ( .A1(id_pc[6]), .A2(n3), .B1(if_pc[6]), .B2(n2), .Z(n10)
         );
  I2NOR3V1_8TH40 U69 ( .A1(flush_BAR), .A2(stall_ctrl[1]), .B(rst), .ZN(n3) );
endmodule


module inst_decode_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:4] carry;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  AD1V2C_8TH40 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  AD1V2C_8TH40 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), 
        .S(SUM[30]) );
  AD1V2C_8TH40 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), 
        .S(SUM[29]) );
  AD1V2C_8TH40 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), 
        .S(SUM[28]) );
  AD1V2C_8TH40 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), 
        .S(SUM[27]) );
  AD1V2C_8TH40 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), 
        .S(SUM[26]) );
  AD1V2C_8TH40 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), 
        .S(SUM[25]) );
  AD1V2C_8TH40 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), 
        .S(SUM[24]) );
  AD1V2C_8TH40 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), 
        .S(SUM[23]) );
  AD1V2C_8TH40 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), 
        .S(SUM[22]) );
  AD1V2C_8TH40 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), 
        .S(SUM[21]) );
  AD1V2C_8TH40 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), 
        .S(SUM[20]) );
  AD1V2C_8TH40 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), 
        .S(SUM[19]) );
  AD1V2C_8TH40 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), 
        .S(SUM[18]) );
  AD1V2C_8TH40 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), 
        .S(SUM[17]) );
  AD1V2C_8TH40 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), 
        .S(SUM[16]) );
  AD1V2C_8TH40 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), 
        .S(SUM[15]) );
  AD1V2C_8TH40 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), 
        .S(SUM[14]) );
  AD1V2C_8TH40 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), 
        .S(SUM[13]) );
  AD1V2C_8TH40 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), 
        .S(SUM[12]) );
  AD1V2C_8TH40 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), 
        .S(SUM[11]) );
  AD1V2C_8TH40 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S(SUM[10]) );
  AD1V2C_8TH40 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  AD1V2C_8TH40 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  AD1V2C_8TH40 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  AD1V2C_8TH40 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  AD1V2C_8TH40 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  AD1V2C_8TH40 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  AD1V2C_8TH40 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3])
         );
  AND2V2_8TH40 U1 ( .A1(A[2]), .A2(B[2]), .Z(n1) );
  XOR2V2_8TH40 U2 ( .A1(A[2]), .A2(B[2]), .Z(SUM[2]) );
endmodule


module inst_decode_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  XNOR2V2_8TH40 U1 ( .A1(A[31]), .A2(n28), .ZN(SUM[31]) );
  NAND2V2_8TH40 U2 ( .A1(n27), .A2(A[30]), .ZN(n28) );
  INV2_8TH40 U3 ( .I(A[2]), .ZN(SUM[2]) );
  AND2V2_8TH40 U4 ( .A1(A[2]), .A2(A[3]), .Z(n1) );
  AND2V2_8TH40 U5 ( .A1(n1), .A2(A[4]), .Z(n2) );
  AND2V2_8TH40 U6 ( .A1(n2), .A2(A[5]), .Z(n3) );
  AND2V2_8TH40 U7 ( .A1(n3), .A2(A[6]), .Z(n4) );
  AND2V2_8TH40 U8 ( .A1(n4), .A2(A[7]), .Z(n5) );
  AND2V2_8TH40 U9 ( .A1(n5), .A2(A[8]), .Z(n6) );
  AND2V2_8TH40 U10 ( .A1(n6), .A2(A[9]), .Z(n7) );
  AND2V2_8TH40 U11 ( .A1(n7), .A2(A[10]), .Z(n8) );
  AND2V2_8TH40 U12 ( .A1(n8), .A2(A[11]), .Z(n9) );
  AND2V2_8TH40 U13 ( .A1(n9), .A2(A[12]), .Z(n10) );
  AND2V2_8TH40 U14 ( .A1(n10), .A2(A[13]), .Z(n11) );
  AND2V2_8TH40 U15 ( .A1(n11), .A2(A[14]), .Z(n12) );
  AND2V2_8TH40 U16 ( .A1(n12), .A2(A[15]), .Z(n13) );
  AND2V2_8TH40 U17 ( .A1(n13), .A2(A[16]), .Z(n14) );
  AND2V2_8TH40 U18 ( .A1(n14), .A2(A[17]), .Z(n15) );
  AND2V2_8TH40 U19 ( .A1(n15), .A2(A[18]), .Z(n16) );
  AND2V2_8TH40 U20 ( .A1(n16), .A2(A[19]), .Z(n17) );
  AND2V2_8TH40 U21 ( .A1(n17), .A2(A[20]), .Z(n18) );
  AND2V2_8TH40 U22 ( .A1(n18), .A2(A[21]), .Z(n19) );
  AND2V2_8TH40 U23 ( .A1(n19), .A2(A[22]), .Z(n20) );
  AND2V2_8TH40 U24 ( .A1(n20), .A2(A[23]), .Z(n21) );
  AND2V2_8TH40 U25 ( .A1(n21), .A2(A[24]), .Z(n22) );
  AND2V2_8TH40 U26 ( .A1(n22), .A2(A[25]), .Z(n23) );
  AND2V2_8TH40 U27 ( .A1(n23), .A2(A[26]), .Z(n24) );
  AND2V2_8TH40 U28 ( .A1(n24), .A2(A[27]), .Z(n25) );
  AND2V2_8TH40 U29 ( .A1(n25), .A2(A[28]), .Z(n26) );
  AND2V2_8TH40 U30 ( .A1(n26), .A2(A[29]), .Z(n27) );
  XOR2V2_8TH40 U31 ( .A1(n27), .A2(A[30]), .Z(SUM[30]) );
  XOR2V2_8TH40 U32 ( .A1(n26), .A2(A[29]), .Z(SUM[29]) );
  XOR2V2_8TH40 U33 ( .A1(n25), .A2(A[28]), .Z(SUM[28]) );
  XOR2V2_8TH40 U34 ( .A1(n24), .A2(A[27]), .Z(SUM[27]) );
  XOR2V2_8TH40 U35 ( .A1(n23), .A2(A[26]), .Z(SUM[26]) );
  XOR2V2_8TH40 U36 ( .A1(n22), .A2(A[25]), .Z(SUM[25]) );
  XOR2V2_8TH40 U37 ( .A1(n21), .A2(A[24]), .Z(SUM[24]) );
  XOR2V2_8TH40 U38 ( .A1(n20), .A2(A[23]), .Z(SUM[23]) );
  XOR2V2_8TH40 U39 ( .A1(n19), .A2(A[22]), .Z(SUM[22]) );
  XOR2V2_8TH40 U40 ( .A1(n18), .A2(A[21]), .Z(SUM[21]) );
  XOR2V2_8TH40 U41 ( .A1(n17), .A2(A[20]), .Z(SUM[20]) );
  XOR2V2_8TH40 U42 ( .A1(n16), .A2(A[19]), .Z(SUM[19]) );
  XOR2V2_8TH40 U43 ( .A1(n15), .A2(A[18]), .Z(SUM[18]) );
  XOR2V2_8TH40 U44 ( .A1(n14), .A2(A[17]), .Z(SUM[17]) );
  XOR2V2_8TH40 U45 ( .A1(n13), .A2(A[16]), .Z(SUM[16]) );
  XOR2V2_8TH40 U46 ( .A1(n12), .A2(A[15]), .Z(SUM[15]) );
  XOR2V2_8TH40 U47 ( .A1(n11), .A2(A[14]), .Z(SUM[14]) );
  XOR2V2_8TH40 U48 ( .A1(n10), .A2(A[13]), .Z(SUM[13]) );
  XOR2V2_8TH40 U49 ( .A1(n9), .A2(A[12]), .Z(SUM[12]) );
  XOR2V2_8TH40 U50 ( .A1(n8), .A2(A[11]), .Z(SUM[11]) );
  XOR2V2_8TH40 U51 ( .A1(n7), .A2(A[10]), .Z(SUM[10]) );
  XOR2V2_8TH40 U52 ( .A1(n6), .A2(A[9]), .Z(SUM[9]) );
  XOR2V2_8TH40 U53 ( .A1(n5), .A2(A[8]), .Z(SUM[8]) );
  XOR2V2_8TH40 U54 ( .A1(n4), .A2(A[7]), .Z(SUM[7]) );
  XOR2V2_8TH40 U55 ( .A1(n3), .A2(A[6]), .Z(SUM[6]) );
  XOR2V2_8TH40 U56 ( .A1(n2), .A2(A[5]), .Z(SUM[5]) );
  XOR2V2_8TH40 U57 ( .A1(n1), .A2(A[4]), .Z(SUM[4]) );
  XOR2V2_8TH40 U58 ( .A1(A[2]), .A2(A[3]), .Z(SUM[3]) );
endmodule


module inst_decode_DW01_cmp6_3 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  AND2V4_8TH40 U1 ( .A1(n4), .A2(n5), .Z(EQ) );
  NOR4V2_8TH40 U2 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  NAND4V2_8TH40 U3 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .ZN(n7) );
  NAND4V2_8TH40 U4 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(n8) );
  NAND4V2_8TH40 U5 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(n9) );
  NOR4V2_8TH40 U6 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NAND4V2_8TH40 U7 ( .A1(n22), .A2(n23), .A3(n24), .A4(n25), .ZN(n6) );
  OAI22V2_8TH40 U8 ( .A1(n26), .A2(n2), .B1(B[1]), .B2(n26), .ZN(n25) );
  NAND4V2_8TH40 U9 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  NAND4V2_8TH40 U10 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  NAND4V2_8TH40 U11 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  NAND4V2_8TH40 U12 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  INV2_8TH40 U13 ( .I(B[1]), .ZN(n3) );
  INV2_8TH40 U14 ( .I(A[1]), .ZN(n2) );
  XNOR2V0_8TH40 U15 ( .A1(B[11]), .A2(A[11]), .ZN(n13) );
  XNOR2V0_8TH40 U16 ( .A1(B[12]), .A2(A[12]), .ZN(n12) );
  XNOR2V0_8TH40 U17 ( .A1(B[13]), .A2(A[13]), .ZN(n11) );
  XNOR2V0_8TH40 U18 ( .A1(B[14]), .A2(A[14]), .ZN(n10) );
  XNOR2V0_8TH40 U19 ( .A1(B[7]), .A2(A[7]), .ZN(n17) );
  XNOR2V0_8TH40 U20 ( .A1(B[8]), .A2(A[8]), .ZN(n16) );
  XNOR2V0_8TH40 U21 ( .A1(B[9]), .A2(A[9]), .ZN(n15) );
  XNOR2V0_8TH40 U22 ( .A1(B[10]), .A2(A[10]), .ZN(n14) );
  XNOR2V0_8TH40 U23 ( .A1(B[3]), .A2(A[3]), .ZN(n21) );
  XNOR2V0_8TH40 U24 ( .A1(B[4]), .A2(A[4]), .ZN(n20) );
  XNOR2V0_8TH40 U25 ( .A1(B[5]), .A2(A[5]), .ZN(n19) );
  XNOR2V0_8TH40 U26 ( .A1(B[6]), .A2(A[6]), .ZN(n18) );
  INOR2V0_8TH40 U27 ( .A1(B[0]), .B1(A[0]), .ZN(n26) );
  OAI22V0_8TH40 U28 ( .A1(A[1]), .A2(n27), .B1(n27), .B2(n3), .ZN(n24) );
  INOR2V0_8TH40 U29 ( .A1(A[0]), .B1(B[0]), .ZN(n27) );
  XNOR2V0_8TH40 U30 ( .A1(B[31]), .A2(A[31]), .ZN(n23) );
  XNOR2V0_8TH40 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n22) );
  XNOR2V0_8TH40 U32 ( .A1(B[27]), .A2(A[27]), .ZN(n35) );
  XNOR2V0_8TH40 U33 ( .A1(B[28]), .A2(A[28]), .ZN(n34) );
  XNOR2V0_8TH40 U34 ( .A1(B[29]), .A2(A[29]), .ZN(n33) );
  XNOR2V0_8TH40 U35 ( .A1(B[30]), .A2(A[30]), .ZN(n32) );
  XNOR2V0_8TH40 U36 ( .A1(B[23]), .A2(A[23]), .ZN(n39) );
  XNOR2V0_8TH40 U37 ( .A1(B[24]), .A2(A[24]), .ZN(n38) );
  XNOR2V0_8TH40 U38 ( .A1(B[25]), .A2(A[25]), .ZN(n37) );
  XNOR2V0_8TH40 U39 ( .A1(B[26]), .A2(A[26]), .ZN(n36) );
  XNOR2V0_8TH40 U40 ( .A1(B[19]), .A2(A[19]), .ZN(n43) );
  XNOR2V0_8TH40 U41 ( .A1(B[20]), .A2(A[20]), .ZN(n42) );
  XNOR2V0_8TH40 U42 ( .A1(B[21]), .A2(A[21]), .ZN(n41) );
  XNOR2V0_8TH40 U43 ( .A1(B[22]), .A2(A[22]), .ZN(n40) );
  XNOR2V0_8TH40 U44 ( .A1(B[15]), .A2(A[15]), .ZN(n47) );
  XNOR2V0_8TH40 U45 ( .A1(B[16]), .A2(A[16]), .ZN(n46) );
  XNOR2V0_8TH40 U46 ( .A1(B[17]), .A2(A[17]), .ZN(n45) );
  XNOR2V0_8TH40 U47 ( .A1(B[18]), .A2(A[18]), .ZN(n44) );
endmodule


module inst_decode_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV2_8TH40 U1 ( .I(A[3]), .ZN(SUM[3]) );
  XNOR2V2_8TH40 U2 ( .A1(A[31]), .A2(n27), .ZN(SUM[31]) );
  NAND2V2_8TH40 U3 ( .A1(n26), .A2(A[30]), .ZN(n27) );
  AND2V2_8TH40 U4 ( .A1(A[3]), .A2(A[4]), .Z(n1) );
  AND2V2_8TH40 U5 ( .A1(n1), .A2(A[5]), .Z(n2) );
  AND2V2_8TH40 U6 ( .A1(n2), .A2(A[6]), .Z(n3) );
  AND2V2_8TH40 U7 ( .A1(n3), .A2(A[7]), .Z(n4) );
  AND2V2_8TH40 U8 ( .A1(n4), .A2(A[8]), .Z(n5) );
  AND2V2_8TH40 U9 ( .A1(n5), .A2(A[9]), .Z(n6) );
  AND2V2_8TH40 U10 ( .A1(n6), .A2(A[10]), .Z(n7) );
  AND2V2_8TH40 U11 ( .A1(n7), .A2(A[11]), .Z(n8) );
  AND2V2_8TH40 U12 ( .A1(n8), .A2(A[12]), .Z(n9) );
  AND2V2_8TH40 U13 ( .A1(n9), .A2(A[13]), .Z(n10) );
  AND2V2_8TH40 U14 ( .A1(n10), .A2(A[14]), .Z(n11) );
  AND2V2_8TH40 U15 ( .A1(n11), .A2(A[15]), .Z(n12) );
  AND2V2_8TH40 U16 ( .A1(n12), .A2(A[16]), .Z(n13) );
  AND2V2_8TH40 U17 ( .A1(n13), .A2(A[17]), .Z(n14) );
  AND2V2_8TH40 U18 ( .A1(n14), .A2(A[18]), .Z(n15) );
  AND2V2_8TH40 U19 ( .A1(n15), .A2(A[19]), .Z(n16) );
  AND2V2_8TH40 U20 ( .A1(n16), .A2(A[20]), .Z(n17) );
  AND2V2_8TH40 U21 ( .A1(n17), .A2(A[21]), .Z(n18) );
  AND2V2_8TH40 U22 ( .A1(n18), .A2(A[22]), .Z(n19) );
  AND2V2_8TH40 U23 ( .A1(n19), .A2(A[23]), .Z(n20) );
  AND2V2_8TH40 U24 ( .A1(n20), .A2(A[24]), .Z(n21) );
  AND2V2_8TH40 U25 ( .A1(n21), .A2(A[25]), .Z(n22) );
  AND2V2_8TH40 U26 ( .A1(n22), .A2(A[26]), .Z(n23) );
  AND2V2_8TH40 U27 ( .A1(n23), .A2(A[27]), .Z(n24) );
  AND2V2_8TH40 U28 ( .A1(n24), .A2(A[28]), .Z(n25) );
  AND2V2_8TH40 U29 ( .A1(n25), .A2(A[29]), .Z(n26) );
  XOR2V2_8TH40 U30 ( .A1(n26), .A2(A[30]), .Z(SUM[30]) );
  XOR2V2_8TH40 U31 ( .A1(n25), .A2(A[29]), .Z(SUM[29]) );
  XOR2V2_8TH40 U32 ( .A1(n24), .A2(A[28]), .Z(SUM[28]) );
  XOR2V2_8TH40 U33 ( .A1(n23), .A2(A[27]), .Z(SUM[27]) );
  XOR2V2_8TH40 U34 ( .A1(n22), .A2(A[26]), .Z(SUM[26]) );
  XOR2V2_8TH40 U35 ( .A1(n21), .A2(A[25]), .Z(SUM[25]) );
  XOR2V2_8TH40 U36 ( .A1(n20), .A2(A[24]), .Z(SUM[24]) );
  XOR2V2_8TH40 U37 ( .A1(n19), .A2(A[23]), .Z(SUM[23]) );
  XOR2V2_8TH40 U38 ( .A1(n18), .A2(A[22]), .Z(SUM[22]) );
  XOR2V2_8TH40 U39 ( .A1(n17), .A2(A[21]), .Z(SUM[21]) );
  XOR2V2_8TH40 U40 ( .A1(n16), .A2(A[20]), .Z(SUM[20]) );
  XOR2V2_8TH40 U41 ( .A1(n15), .A2(A[19]), .Z(SUM[19]) );
  XOR2V2_8TH40 U42 ( .A1(n14), .A2(A[18]), .Z(SUM[18]) );
  XOR2V2_8TH40 U43 ( .A1(n13), .A2(A[17]), .Z(SUM[17]) );
  XOR2V2_8TH40 U44 ( .A1(n12), .A2(A[16]), .Z(SUM[16]) );
  XOR2V2_8TH40 U45 ( .A1(n11), .A2(A[15]), .Z(SUM[15]) );
  XOR2V2_8TH40 U46 ( .A1(n10), .A2(A[14]), .Z(SUM[14]) );
  XOR2V2_8TH40 U47 ( .A1(n9), .A2(A[13]), .Z(SUM[13]) );
  XOR2V2_8TH40 U48 ( .A1(n8), .A2(A[12]), .Z(SUM[12]) );
  XOR2V2_8TH40 U49 ( .A1(n7), .A2(A[11]), .Z(SUM[11]) );
  XOR2V2_8TH40 U50 ( .A1(n6), .A2(A[10]), .Z(SUM[10]) );
  XOR2V2_8TH40 U51 ( .A1(n5), .A2(A[9]), .Z(SUM[9]) );
  XOR2V2_8TH40 U52 ( .A1(n4), .A2(A[8]), .Z(SUM[8]) );
  XOR2V2_8TH40 U53 ( .A1(n3), .A2(A[7]), .Z(SUM[7]) );
  XOR2V2_8TH40 U54 ( .A1(n2), .A2(A[6]), .Z(SUM[6]) );
  XOR2V2_8TH40 U55 ( .A1(n1), .A2(A[5]), .Z(SUM[5]) );
  XOR2V2_8TH40 U56 ( .A1(A[3]), .A2(A[4]), .Z(SUM[4]) );
endmodule


module inst_decode ( rst, pc_i, inst_i, gpr1_data_i, gpr2_data_i, 
        df_exid_gpr_we, df_exid_target_gpr, df_exid_exe_result, 
        df_memid_gpr_we, df_memid_target_gpr, df_memid_exe_result, 
        curid_inst_delayslot_i, ex_inst_type, gpr1_re, gpr2_re, gpr1_addr, 
        gpr2_addr, inst_type, inst_class, gpr1_data_o, gpr2_data_o, target_gpr, 
        gpr_we, stall_req, branch_flag, branch_target_addr, link_addr, 
        nxtid_inst_delayslot_o, curid_inst_delayslot_o, inst_o, except_type, 
        cur_inst_addr );
  input [31:0] pc_i;
  input [31:0] inst_i;
  input [31:0] gpr1_data_i;
  input [31:0] gpr2_data_i;
  input [4:0] df_exid_target_gpr;
  input [31:0] df_exid_exe_result;
  input [4:0] df_memid_target_gpr;
  input [31:0] df_memid_exe_result;
  input [7:0] ex_inst_type;
  output [4:0] gpr1_addr;
  output [4:0] gpr2_addr;
  output [7:0] inst_type;
  output [2:0] inst_class;
  output [31:0] gpr1_data_o;
  output [31:0] gpr2_data_o;
  output [4:0] target_gpr;
  output [31:0] branch_target_addr;
  output [31:0] link_addr;
  output [31:0] inst_o;
  output [31:0] except_type;
  output [31:0] cur_inst_addr;
  input rst, df_exid_gpr_we, df_memid_gpr_we, curid_inst_delayslot_i;
  output gpr1_re, gpr2_re, gpr_we, stall_req, branch_flag,
         nxtid_inst_delayslot_o, curid_inst_delayslot_o;
  wire   branch_flag, N812, N1698, N1699, N1700, N1701, N1702, N1703, N1704,
         N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714,
         N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724,
         N1725, N1726, N1727, N1728, N1729, N1730, N1756, N1757, N1758, N1759,
         N1760, N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, N1769,
         N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779,
         N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n1, n2, n3, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507;
  wire   [31:0] pc_plus8;
  wire   [31:0] pc_plus4;
  assign nxtid_inst_delayslot_o = branch_flag;
  assign inst_o[15] = inst_i[15];
  assign inst_o[14] = inst_i[14];
  assign inst_o[13] = inst_i[13];
  assign inst_o[12] = inst_i[12];
  assign inst_o[11] = inst_i[11];
  assign inst_o[10] = inst_i[10];
  assign inst_o[9] = inst_i[9];
  assign inst_o[8] = inst_i[8];
  assign inst_o[7] = inst_i[7];
  assign inst_o[6] = inst_i[6];
  assign inst_o[5] = inst_i[5];
  assign inst_o[4] = inst_i[4];
  assign inst_o[3] = inst_i[3];
  assign inst_o[2] = inst_i[2];
  assign inst_o[1] = inst_i[1];
  assign inst_o[0] = inst_i[0];
  assign cur_inst_addr[31] = pc_i[31];
  assign cur_inst_addr[30] = pc_i[30];
  assign cur_inst_addr[29] = pc_i[29];
  assign cur_inst_addr[28] = pc_i[28];
  assign cur_inst_addr[27] = pc_i[27];
  assign cur_inst_addr[26] = pc_i[26];
  assign cur_inst_addr[25] = pc_i[25];
  assign cur_inst_addr[24] = pc_i[24];
  assign cur_inst_addr[23] = pc_i[23];
  assign cur_inst_addr[22] = pc_i[22];
  assign cur_inst_addr[21] = pc_i[21];
  assign cur_inst_addr[20] = pc_i[20];
  assign cur_inst_addr[19] = pc_i[19];
  assign cur_inst_addr[18] = pc_i[18];
  assign cur_inst_addr[17] = pc_i[17];
  assign cur_inst_addr[16] = pc_i[16];
  assign cur_inst_addr[15] = pc_i[15];
  assign cur_inst_addr[14] = pc_i[14];
  assign cur_inst_addr[13] = pc_i[13];
  assign cur_inst_addr[12] = pc_i[12];
  assign cur_inst_addr[11] = pc_i[11];
  assign cur_inst_addr[10] = pc_i[10];
  assign cur_inst_addr[9] = pc_i[9];
  assign cur_inst_addr[8] = pc_i[8];
  assign cur_inst_addr[7] = pc_i[7];
  assign cur_inst_addr[6] = pc_i[6];
  assign cur_inst_addr[5] = pc_i[5];
  assign cur_inst_addr[4] = pc_i[4];
  assign cur_inst_addr[3] = pc_i[3];
  assign cur_inst_addr[2] = pc_i[2];
  assign cur_inst_addr[1] = pc_i[1];
  assign cur_inst_addr[0] = pc_i[0];

  LAHQV1_8TH40 gpr1_data_o_reg_31_ ( .E(N1698), .D(N1730), .Q(gpr1_data_o[31])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_30_ ( .E(N1698), .D(N1729), .Q(gpr1_data_o[30])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_29_ ( .E(N1698), .D(N1728), .Q(gpr1_data_o[29])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_28_ ( .E(N1698), .D(N1727), .Q(gpr1_data_o[28])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_27_ ( .E(N1698), .D(N1726), .Q(gpr1_data_o[27])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_26_ ( .E(N1698), .D(N1725), .Q(gpr1_data_o[26])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_25_ ( .E(N1698), .D(N1724), .Q(gpr1_data_o[25])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_24_ ( .E(N1698), .D(N1723), .Q(gpr1_data_o[24])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_23_ ( .E(N1698), .D(N1722), .Q(gpr1_data_o[23])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_22_ ( .E(N1698), .D(N1721), .Q(gpr1_data_o[22])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_21_ ( .E(N1698), .D(N1720), .Q(gpr1_data_o[21])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_20_ ( .E(N1698), .D(N1719), .Q(gpr1_data_o[20])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_19_ ( .E(N1698), .D(N1718), .Q(gpr1_data_o[19])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_18_ ( .E(N1698), .D(N1717), .Q(gpr1_data_o[18])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_17_ ( .E(N1698), .D(N1716), .Q(gpr1_data_o[17])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_16_ ( .E(N1698), .D(N1715), .Q(gpr1_data_o[16])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_15_ ( .E(N1698), .D(N1714), .Q(gpr1_data_o[15])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_14_ ( .E(N1698), .D(N1713), .Q(gpr1_data_o[14])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_13_ ( .E(N1698), .D(N1712), .Q(gpr1_data_o[13])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_12_ ( .E(N1698), .D(N1711), .Q(gpr1_data_o[12])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_11_ ( .E(N1698), .D(N1710), .Q(gpr1_data_o[11])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_10_ ( .E(N1698), .D(N1709), .Q(gpr1_data_o[10])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_9_ ( .E(N1698), .D(N1708), .Q(gpr1_data_o[9])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_8_ ( .E(N1698), .D(N1707), .Q(gpr1_data_o[8])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_7_ ( .E(N1698), .D(N1706), .Q(gpr1_data_o[7])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_6_ ( .E(N1698), .D(N1705), .Q(gpr1_data_o[6])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_5_ ( .E(N1698), .D(N1704), .Q(gpr1_data_o[5])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_4_ ( .E(N1698), .D(N1703), .Q(gpr1_data_o[4])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_3_ ( .E(N1698), .D(N1702), .Q(gpr1_data_o[3])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_2_ ( .E(N1698), .D(N1701), .Q(gpr1_data_o[2])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_1_ ( .E(N1698), .D(N1700), .Q(gpr1_data_o[1])
         );
  LAHQV1_8TH40 gpr1_data_o_reg_0_ ( .E(N1698), .D(N1699), .Q(gpr1_data_o[0])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_31_ ( .E(N1756), .D(N1788), .Q(gpr2_data_o[31])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_30_ ( .E(N1756), .D(N1787), .Q(gpr2_data_o[30])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_29_ ( .E(N1756), .D(N1786), .Q(gpr2_data_o[29])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_28_ ( .E(N1756), .D(N1785), .Q(gpr2_data_o[28])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_27_ ( .E(N1756), .D(N1784), .Q(gpr2_data_o[27])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_26_ ( .E(N1756), .D(N1783), .Q(gpr2_data_o[26])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_25_ ( .E(N1756), .D(N1782), .Q(gpr2_data_o[25])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_24_ ( .E(N1756), .D(N1781), .Q(gpr2_data_o[24])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_23_ ( .E(N1756), .D(N1780), .Q(gpr2_data_o[23])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_22_ ( .E(N1756), .D(N1779), .Q(gpr2_data_o[22])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_21_ ( .E(N1756), .D(N1778), .Q(gpr2_data_o[21])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_20_ ( .E(N1756), .D(N1777), .Q(gpr2_data_o[20])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_19_ ( .E(N1756), .D(N1776), .Q(gpr2_data_o[19])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_18_ ( .E(N1756), .D(N1775), .Q(gpr2_data_o[18])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_17_ ( .E(N1756), .D(N1774), .Q(gpr2_data_o[17])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_16_ ( .E(N1756), .D(N1773), .Q(gpr2_data_o[16])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_15_ ( .E(N1756), .D(N1772), .Q(gpr2_data_o[15])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_14_ ( .E(N1756), .D(N1771), .Q(gpr2_data_o[14])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_13_ ( .E(N1756), .D(N1770), .Q(gpr2_data_o[13])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_12_ ( .E(N1756), .D(N1769), .Q(gpr2_data_o[12])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_11_ ( .E(N1756), .D(N1768), .Q(gpr2_data_o[11])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_10_ ( .E(N1756), .D(N1767), .Q(gpr2_data_o[10])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_9_ ( .E(N1756), .D(N1766), .Q(gpr2_data_o[9])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_8_ ( .E(N1756), .D(N1765), .Q(gpr2_data_o[8])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_7_ ( .E(N1756), .D(N1764), .Q(gpr2_data_o[7])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_6_ ( .E(N1756), .D(N1763), .Q(gpr2_data_o[6])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_5_ ( .E(N1756), .D(N1762), .Q(gpr2_data_o[5])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_4_ ( .E(N1756), .D(N1761), .Q(gpr2_data_o[4])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_3_ ( .E(N1756), .D(N1760), .Q(gpr2_data_o[3])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_2_ ( .E(N1756), .D(N1759), .Q(gpr2_data_o[2])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_1_ ( .E(N1756), .D(N1758), .Q(gpr2_data_o[1])
         );
  LAHQV1_8TH40 gpr2_data_o_reg_0_ ( .E(N1756), .D(N1757), .Q(gpr2_data_o[0])
         );
  inst_decode_DW01_add_0 r221 ( .A(pc_plus4), .B({inst_i[15], inst_i[15], 
        inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], 
        inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], 
        inst_i[15:0], 1'b0, 1'b0}), .CI(1'b0), .SUM({n4, n5, n6, n7, n8, n9, 
        n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
        n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35}) );
  inst_decode_DW01_add_1 add_76 ( .A(pc_i), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(pc_plus4) );
  inst_decode_DW01_cmp6_3 r238 ( .A(gpr1_data_o), .B(gpr2_data_o), .TC(1'b0), 
        .EQ(N812) );
  inst_decode_DW01_add_2 add_75 ( .A(pc_i), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(pc_plus8) );
  NOR3V2_8TH40 U3 ( .A1(n444), .A2(n446), .A3(n445), .ZN(n399) );
  AO222V4_8TH40 U4 ( .A1(n399), .A2(df_exid_exe_result[31]), .B1(n400), .B2(
        df_memid_exe_result[31]), .C1(gpr1_data_i[31]), .C2(n401), .Z(N1730)
         );
  AO222V4_8TH40 U5 ( .A1(n399), .A2(df_exid_exe_result[30]), .B1(n400), .B2(
        df_memid_exe_result[30]), .C1(gpr1_data_i[30]), .C2(n401), .Z(N1729)
         );
  AO222V4_8TH40 U6 ( .A1(n399), .A2(df_exid_exe_result[29]), .B1(n400), .B2(
        df_memid_exe_result[29]), .C1(gpr1_data_i[29]), .C2(n401), .Z(N1728)
         );
  AO222V4_8TH40 U7 ( .A1(n399), .A2(df_exid_exe_result[28]), .B1(n400), .B2(
        df_memid_exe_result[28]), .C1(gpr1_data_i[28]), .C2(n401), .Z(N1727)
         );
  AO222V4_8TH40 U8 ( .A1(n399), .A2(df_exid_exe_result[27]), .B1(n400), .B2(
        df_memid_exe_result[27]), .C1(gpr1_data_i[27]), .C2(n401), .Z(N1726)
         );
  AO222V4_8TH40 U9 ( .A1(n399), .A2(df_exid_exe_result[26]), .B1(n400), .B2(
        df_memid_exe_result[26]), .C1(gpr1_data_i[26]), .C2(n401), .Z(N1725)
         );
  AO222V4_8TH40 U10 ( .A1(n399), .A2(df_exid_exe_result[25]), .B1(n400), .B2(
        df_memid_exe_result[25]), .C1(gpr1_data_i[25]), .C2(n401), .Z(N1724)
         );
  AO222V4_8TH40 U11 ( .A1(n399), .A2(df_exid_exe_result[24]), .B1(n400), .B2(
        df_memid_exe_result[24]), .C1(gpr1_data_i[24]), .C2(n401), .Z(N1723)
         );
  AO222V4_8TH40 U12 ( .A1(n399), .A2(df_exid_exe_result[23]), .B1(n400), .B2(
        df_memid_exe_result[23]), .C1(gpr1_data_i[23]), .C2(n401), .Z(N1722)
         );
  AO222V4_8TH40 U13 ( .A1(n399), .A2(df_exid_exe_result[22]), .B1(n400), .B2(
        df_memid_exe_result[22]), .C1(gpr1_data_i[22]), .C2(n401), .Z(N1721)
         );
  AO222V4_8TH40 U14 ( .A1(n399), .A2(df_exid_exe_result[21]), .B1(n400), .B2(
        df_memid_exe_result[21]), .C1(gpr1_data_i[21]), .C2(n401), .Z(N1720)
         );
  AO222V4_8TH40 U15 ( .A1(n399), .A2(df_exid_exe_result[20]), .B1(n400), .B2(
        df_memid_exe_result[20]), .C1(gpr1_data_i[20]), .C2(n401), .Z(N1719)
         );
  AO222V4_8TH40 U16 ( .A1(n399), .A2(df_exid_exe_result[19]), .B1(n400), .B2(
        df_memid_exe_result[19]), .C1(gpr1_data_i[19]), .C2(n401), .Z(N1718)
         );
  AO222V4_8TH40 U17 ( .A1(n399), .A2(df_exid_exe_result[18]), .B1(n400), .B2(
        df_memid_exe_result[18]), .C1(gpr1_data_i[18]), .C2(n401), .Z(N1717)
         );
  AO222V4_8TH40 U18 ( .A1(n399), .A2(df_exid_exe_result[17]), .B1(n400), .B2(
        df_memid_exe_result[17]), .C1(gpr1_data_i[17]), .C2(n401), .Z(N1716)
         );
  AO222V4_8TH40 U19 ( .A1(n399), .A2(df_exid_exe_result[16]), .B1(n400), .B2(
        df_memid_exe_result[16]), .C1(gpr1_data_i[16]), .C2(n401), .Z(N1715)
         );
  OAI31V2_8TH40 U20 ( .A1(n467), .A2(n181), .A3(n164), .B(n468), .ZN(n466) );
  INOR2V4_8TH40 U21 ( .A1(pc_plus8[5]), .B1(n59), .ZN(link_addr[5]) );
  INOR2V4_8TH40 U22 ( .A1(pc_plus8[6]), .B1(n59), .ZN(link_addr[6]) );
  INOR2V4_8TH40 U23 ( .A1(pc_plus8[7]), .B1(n59), .ZN(link_addr[7]) );
  INOR2V4_8TH40 U24 ( .A1(pc_plus8[8]), .B1(n59), .ZN(link_addr[8]) );
  INOR2V4_8TH40 U25 ( .A1(pc_plus8[9]), .B1(n59), .ZN(link_addr[9]) );
  INOR2V4_8TH40 U26 ( .A1(pc_plus8[10]), .B1(n59), .ZN(link_addr[10]) );
  INOR2V4_8TH40 U27 ( .A1(pc_plus8[11]), .B1(n59), .ZN(link_addr[11]) );
  INOR2V4_8TH40 U28 ( .A1(pc_plus8[12]), .B1(n59), .ZN(link_addr[12]) );
  INOR2V4_8TH40 U29 ( .A1(pc_plus8[13]), .B1(n59), .ZN(link_addr[13]) );
  INOR2V4_8TH40 U30 ( .A1(pc_plus8[14]), .B1(n59), .ZN(link_addr[14]) );
  INOR2V4_8TH40 U31 ( .A1(pc_plus8[15]), .B1(n59), .ZN(link_addr[15]) );
  INOR2V4_8TH40 U32 ( .A1(pc_plus8[16]), .B1(n59), .ZN(link_addr[16]) );
  INOR2V4_8TH40 U33 ( .A1(pc_plus8[17]), .B1(n59), .ZN(link_addr[17]) );
  INOR2V4_8TH40 U34 ( .A1(pc_plus8[18]), .B1(n59), .ZN(link_addr[18]) );
  INOR2V4_8TH40 U35 ( .A1(pc_plus8[19]), .B1(n59), .ZN(link_addr[19]) );
  INOR2V4_8TH40 U36 ( .A1(pc_plus8[20]), .B1(n59), .ZN(link_addr[20]) );
  INOR2V4_8TH40 U37 ( .A1(pc_plus8[21]), .B1(n59), .ZN(link_addr[21]) );
  INOR2V4_8TH40 U38 ( .A1(pc_plus8[22]), .B1(n59), .ZN(link_addr[22]) );
  INOR2V4_8TH40 U39 ( .A1(pc_plus8[23]), .B1(n59), .ZN(link_addr[23]) );
  INOR2V4_8TH40 U40 ( .A1(pc_plus8[24]), .B1(n59), .ZN(link_addr[24]) );
  INOR2V4_8TH40 U41 ( .A1(pc_plus8[25]), .B1(n59), .ZN(link_addr[25]) );
  INOR2V4_8TH40 U42 ( .A1(pc_plus8[26]), .B1(n59), .ZN(link_addr[26]) );
  INOR2V4_8TH40 U43 ( .A1(pc_plus8[27]), .B1(n59), .ZN(link_addr[27]) );
  INOR2V4_8TH40 U44 ( .A1(pc_plus8[28]), .B1(n59), .ZN(link_addr[28]) );
  INOR2V4_8TH40 U45 ( .A1(pc_plus8[29]), .B1(n59), .ZN(link_addr[29]) );
  INOR2V4_8TH40 U46 ( .A1(pc_plus8[30]), .B1(n59), .ZN(link_addr[30]) );
  INOR2V4_8TH40 U47 ( .A1(pc_plus8[4]), .B1(n59), .ZN(link_addr[4]) );
  MUX2NV2_8TH40 U48 ( .I0(n481), .I1(n482), .S(ex_inst_type[4]), .ZN(n480) );
  INOR2V4_8TH40 U49 ( .A1(pc_plus8[31]), .B1(n59), .ZN(link_addr[31]) );
  INOR2V4_8TH40 U50 ( .A1(pc_plus8[3]), .B1(n59), .ZN(link_addr[3]) );
  CLKNV4_8TH40 U51 ( .I(n43), .ZN(gpr2_addr[3]) );
  NAND2V0_8TH40 U52 ( .A1(inst_i[19]), .A2(n51), .ZN(n43) );
  AO22V4_8TH40 U53 ( .A1(n489), .A2(inst_i[24]), .B1(gpr2_addr[3]), .B2(n71), 
        .Z(gpr1_addr[3]) );
  AOI21V4_8TH40 U54 ( .A1(n45), .A2(n490), .B(n473), .ZN(gpr1_addr[2]) );
  XOR2V0_8TH40 U55 ( .A1(df_memid_target_gpr[3]), .A2(gpr2_addr[3]), .Z(n381)
         );
  OAI211V2_8TH40 U56 ( .A1(n212), .A2(n213), .B(n214), .C(n199), .ZN(n207) );
  I2NOR3V2_8TH40 U57 ( .A1(n161), .A2(n474), .B(n70), .ZN(n248) );
  INV2_8TH40 U58 ( .I(n45), .ZN(gpr2_addr[2]) );
  NAND2V2_8TH40 U59 ( .A1(n51), .A2(n220), .ZN(n59) );
  OAI31V2_8TH40 U60 ( .A1(n221), .A2(n177), .A3(n87), .B(n50), .ZN(n220) );
  OAOI211V2_8TH40 U61 ( .A1(n183), .A2(n478), .B(n182), .C(n129), .ZN(n239) );
  OAI31V2_8TH40 U62 ( .A1(n461), .A2(n71), .A3(n95), .B(n51), .ZN(n445) );
  OAI221V2_8TH40 U63 ( .A1(n180), .A2(n333), .B1(n278), .B2(n373), .C(n374), 
        .ZN(N1757) );
  AOI22V2_8TH40 U64 ( .A1(gpr2_data_i[0]), .A2(n281), .B1(
        df_memid_exe_result[0]), .B2(n332), .ZN(n374) );
  OAI221V2_8TH40 U65 ( .A1(n370), .A2(n333), .B1(n278), .B2(n371), .C(n372), 
        .ZN(N1758) );
  AOI22V2_8TH40 U66 ( .A1(gpr2_data_i[1]), .A2(n281), .B1(
        df_memid_exe_result[1]), .B2(n332), .ZN(n372) );
  OAI221V2_8TH40 U67 ( .A1(n367), .A2(n333), .B1(n278), .B2(n368), .C(n369), 
        .ZN(N1759) );
  AOI22V2_8TH40 U68 ( .A1(gpr2_data_i[2]), .A2(n281), .B1(
        df_memid_exe_result[2]), .B2(n332), .ZN(n369) );
  OAI221V2_8TH40 U69 ( .A1(n364), .A2(n333), .B1(n278), .B2(n365), .C(n366), 
        .ZN(N1760) );
  AOI22V2_8TH40 U70 ( .A1(gpr2_data_i[3]), .A2(n281), .B1(
        df_memid_exe_result[3]), .B2(n332), .ZN(n366) );
  OAI221V2_8TH40 U71 ( .A1(n361), .A2(n333), .B1(n278), .B2(n362), .C(n363), 
        .ZN(N1761) );
  AOI22V2_8TH40 U72 ( .A1(gpr2_data_i[4]), .A2(n281), .B1(
        df_memid_exe_result[4]), .B2(n332), .ZN(n363) );
  OAI221V2_8TH40 U73 ( .A1(n158), .A2(n333), .B1(n278), .B2(n359), .C(n360), 
        .ZN(N1762) );
  AOI22V2_8TH40 U74 ( .A1(gpr2_data_i[5]), .A2(n281), .B1(
        df_memid_exe_result[5]), .B2(n332), .ZN(n360) );
  OAI221V2_8TH40 U75 ( .A1(n356), .A2(n333), .B1(n278), .B2(n357), .C(n358), 
        .ZN(N1763) );
  AOI22V2_8TH40 U76 ( .A1(gpr2_data_i[6]), .A2(n281), .B1(
        df_memid_exe_result[6]), .B2(n332), .ZN(n358) );
  OAI221V2_8TH40 U77 ( .A1(n353), .A2(n333), .B1(n278), .B2(n354), .C(n355), 
        .ZN(N1764) );
  AOI22V2_8TH40 U78 ( .A1(gpr2_data_i[7]), .A2(n281), .B1(
        df_memid_exe_result[7]), .B2(n332), .ZN(n355) );
  OAI221V2_8TH40 U79 ( .A1(n350), .A2(n333), .B1(n278), .B2(n351), .C(n352), 
        .ZN(N1765) );
  AOI22V2_8TH40 U80 ( .A1(gpr2_data_i[8]), .A2(n281), .B1(
        df_memid_exe_result[8]), .B2(n332), .ZN(n352) );
  OAI221V2_8TH40 U81 ( .A1(n347), .A2(n333), .B1(n278), .B2(n348), .C(n349), 
        .ZN(N1766) );
  AOI22V2_8TH40 U82 ( .A1(gpr2_data_i[9]), .A2(n281), .B1(
        df_memid_exe_result[9]), .B2(n332), .ZN(n349) );
  OAI221V2_8TH40 U83 ( .A1(n344), .A2(n333), .B1(n278), .B2(n345), .C(n346), 
        .ZN(N1767) );
  AOI22V2_8TH40 U88 ( .A1(gpr2_data_i[10]), .A2(n281), .B1(
        df_memid_exe_result[10]), .B2(n332), .ZN(n346) );
  OAI221V2_8TH40 U89 ( .A1(n48), .A2(n333), .B1(n278), .B2(n342), .C(n343), 
        .ZN(N1768) );
  AOI22V2_8TH40 U90 ( .A1(gpr2_data_i[11]), .A2(n281), .B1(
        df_memid_exe_result[11]), .B2(n332), .ZN(n343) );
  OAI221V2_8TH40 U91 ( .A1(n46), .A2(n333), .B1(n278), .B2(n340), .C(n341), 
        .ZN(N1769) );
  AOI22V2_8TH40 U92 ( .A1(gpr2_data_i[12]), .A2(n281), .B1(
        df_memid_exe_result[12]), .B2(n332), .ZN(n341) );
  OAI221V2_8TH40 U93 ( .A1(n44), .A2(n333), .B1(n278), .B2(n338), .C(n339), 
        .ZN(N1770) );
  AOI22V2_8TH40 U94 ( .A1(gpr2_data_i[13]), .A2(n281), .B1(
        df_memid_exe_result[13]), .B2(n332), .ZN(n339) );
  OAI221V2_8TH40 U95 ( .A1(n42), .A2(n333), .B1(n278), .B2(n336), .C(n337), 
        .ZN(N1771) );
  AOI22V2_8TH40 U96 ( .A1(gpr2_data_i[14]), .A2(n281), .B1(
        df_memid_exe_result[14]), .B2(n332), .ZN(n337) );
  OAI221V2_8TH40 U97 ( .A1(n2), .A2(n333), .B1(n278), .B2(n334), .C(n335), 
        .ZN(N1772) );
  AOI22V2_8TH40 U98 ( .A1(gpr2_data_i[15]), .A2(n281), .B1(
        df_memid_exe_result[15]), .B2(n332), .ZN(n335) );
  OAI31V2_8TH40 U99 ( .A1(n386), .A2(n387), .A3(n388), .B(n51), .ZN(n380) );
  I2NAND3V2_8TH40 U100 ( .A1(n390), .A2(n211), .B(n56), .ZN(n386) );
  OAI22V2_8TH40 U101 ( .A1(n389), .A2(n87), .B1(n239), .B2(n125), .ZN(n388) );
  INOR4V2_8TH40 U102 ( .A1(df_memid_gpr_we), .B1(n380), .B2(n381), .B3(n382), 
        .ZN(n379) );
  AOI211V2_8TH40 U103 ( .A1(n92), .A2(n178), .B(n179), .C(n107), .ZN(n85) );
  INOR4V2_8TH40 U104 ( .A1(n56), .B1(n100), .B2(n101), .B3(n78), .ZN(n99) );
  AOAI211V2_8TH40 U105 ( .A1(n102), .A2(n103), .B(n87), .C(n104), .ZN(n101) );
  I2NOR4V2_8TH40 U106 ( .A1(n463), .A2(n503), .B1(n251), .B2(n81), .ZN(n55) );
  AOI211V2_8TH40 U107 ( .A1(n256), .A2(n213), .B(n504), .C(n505), .ZN(n503) );
  AOI31V2_8TH40 U108 ( .A1(n147), .A2(n191), .A3(n506), .B(n496), .ZN(n505) );
  OAI211V2_8TH40 U109 ( .A1(n160), .A2(n475), .B(n201), .C(n124), .ZN(n70) );
  NOR4V2_8TH40 U110 ( .A1(n156), .A2(n157), .A3(n109), .A4(n90), .ZN(n153) );
  AOI22V2_8TH40 U111 ( .A1(n175), .A2(n467), .B1(n476), .B2(n174), .ZN(n210)
         );
  OAI221V2_8TH40 U112 ( .A1(n158), .A2(n402), .B1(n424), .B2(n404), .C(n425), 
        .ZN(N1704) );
  AOI22V1_8TH40 U113 ( .A1(n399), .A2(df_exid_exe_result[5]), .B1(
        gpr1_data_i[5]), .B2(n401), .ZN(n425) );
  OAI221V2_8TH40 U114 ( .A1(n356), .A2(n402), .B1(n422), .B2(n404), .C(n423), 
        .ZN(N1705) );
  AOI22V2_8TH40 U115 ( .A1(n399), .A2(df_exid_exe_result[6]), .B1(
        gpr1_data_i[6]), .B2(n401), .ZN(n423) );
  OAI221V2_8TH40 U116 ( .A1(n353), .A2(n402), .B1(n420), .B2(n404), .C(n421), 
        .ZN(N1706) );
  AOI22V2_8TH40 U117 ( .A1(n399), .A2(df_exid_exe_result[7]), .B1(
        gpr1_data_i[7]), .B2(n401), .ZN(n421) );
  OAI221V2_8TH40 U118 ( .A1(n350), .A2(n402), .B1(n418), .B2(n404), .C(n419), 
        .ZN(N1707) );
  AOI22V2_8TH40 U119 ( .A1(n399), .A2(df_exid_exe_result[8]), .B1(
        gpr1_data_i[8]), .B2(n401), .ZN(n419) );
  OAI221V2_8TH40 U120 ( .A1(n347), .A2(n402), .B1(n416), .B2(n404), .C(n417), 
        .ZN(N1708) );
  AOI22V2_8TH40 U121 ( .A1(n399), .A2(df_exid_exe_result[9]), .B1(
        gpr1_data_i[9]), .B2(n401), .ZN(n417) );
  OAI221V2_8TH40 U122 ( .A1(n344), .A2(n402), .B1(n414), .B2(n404), .C(n415), 
        .ZN(N1709) );
  AOI22V2_8TH40 U123 ( .A1(n399), .A2(df_exid_exe_result[10]), .B1(
        gpr1_data_i[10]), .B2(n401), .ZN(n415) );
  OAI221V2_8TH40 U124 ( .A1(n48), .A2(n402), .B1(n412), .B2(n404), .C(n413), 
        .ZN(N1710) );
  AOI22V2_8TH40 U125 ( .A1(n399), .A2(df_exid_exe_result[11]), .B1(
        gpr1_data_i[11]), .B2(n401), .ZN(n413) );
  OAI221V2_8TH40 U126 ( .A1(n46), .A2(n402), .B1(n410), .B2(n404), .C(n411), 
        .ZN(N1711) );
  AOI22V2_8TH40 U127 ( .A1(n399), .A2(df_exid_exe_result[12]), .B1(
        gpr1_data_i[12]), .B2(n401), .ZN(n411) );
  OAI221V2_8TH40 U128 ( .A1(n44), .A2(n402), .B1(n408), .B2(n404), .C(n409), 
        .ZN(N1712) );
  AOI22V2_8TH40 U129 ( .A1(n399), .A2(df_exid_exe_result[13]), .B1(
        gpr1_data_i[13]), .B2(n401), .ZN(n409) );
  OAI221V2_8TH40 U130 ( .A1(n42), .A2(n402), .B1(n406), .B2(n404), .C(n407), 
        .ZN(N1713) );
  AOI22V2_8TH40 U131 ( .A1(n399), .A2(df_exid_exe_result[14]), .B1(
        gpr1_data_i[14]), .B2(n401), .ZN(n407) );
  OAI221V2_8TH40 U132 ( .A1(n2), .A2(n402), .B1(n403), .B2(n404), .C(n405), 
        .ZN(N1714) );
  AOI22V2_8TH40 U133 ( .A1(n399), .A2(df_exid_exe_result[15]), .B1(
        gpr1_data_i[15]), .B2(n401), .ZN(n405) );
  OAI211V2_8TH40 U134 ( .A1(n151), .A2(n139), .B(n195), .C(n196), .ZN(n131) );
  I2NOR4V2_8TH40 U135 ( .A1(n118), .A2(n119), .B1(n120), .B2(n78), .ZN(n117)
         );
  INAND4V2_8TH40 U136 ( .A1(n74), .B1(n187), .B2(n188), .B3(n189), .ZN(n137)
         );
  OAI211V2_8TH40 U137 ( .A1(n177), .A2(n224), .B(n201), .C(n225), .ZN(n222) );
  NOR2V2_8TH40 U138 ( .A1(n229), .A2(n230), .ZN(n228) );
  NAND2V2_8TH40 U139 ( .A1(n51), .A2(n52), .ZN(n1) );
  NAND4V2_8TH40 U140 ( .A1(gpr1_re), .A2(df_memid_gpr_we), .A3(n454), .A4(n455), .ZN(n443) );
  NOR4V2_8TH40 U141 ( .A1(n456), .A2(n457), .A3(n458), .A4(n459), .ZN(n455) );
  NAND4V2_8TH40 U142 ( .A1(n376), .A2(n377), .A3(n378), .A4(n379), .ZN(n375)
         );
  I2NOR3V2_8TH40 U143 ( .A1(n192), .A2(n500), .B(n82), .ZN(n242) );
  NAND2V2_8TH40 U144 ( .A1(n51), .A2(n491), .ZN(n490) );
  NAND4V2_8TH40 U145 ( .A1(n119), .A2(n195), .A3(n55), .A4(n492), .ZN(n491) );
  OA211V2_8TH40 U146 ( .A1(n239), .A2(n125), .B(n240), .C(n77), .Z(n203) );
  NAND2V2_8TH40 U147 ( .A1(n470), .A2(n155), .ZN(n112) );
  AOA211V2_8TH40 U148 ( .A1(n169), .A2(n260), .B(n261), .C(n51), .Z(n258) );
  AOI21V2_8TH40 U149 ( .A1(n262), .A2(n263), .B(n264), .ZN(n261) );
  OAI221V2_8TH40 U150 ( .A1(n276), .A2(n326), .B1(n278), .B2(n327), .C(n328), 
        .ZN(N1773) );
  AOI221V2_8TH40 U151 ( .A1(gpr2_data_i[16]), .A2(n281), .B1(n282), .B2(
        inst_i[0]), .C(n283), .ZN(n328) );
  OAI221V2_8TH40 U152 ( .A1(n276), .A2(n323), .B1(n278), .B2(n324), .C(n325), 
        .ZN(N1774) );
  AOI221V2_8TH40 U153 ( .A1(gpr2_data_i[17]), .A2(n281), .B1(n282), .B2(
        inst_i[1]), .C(n283), .ZN(n325) );
  OAI221V2_8TH40 U154 ( .A1(n276), .A2(n320), .B1(n278), .B2(n321), .C(n322), 
        .ZN(N1775) );
  AOI221V2_8TH40 U155 ( .A1(gpr2_data_i[18]), .A2(n281), .B1(n282), .B2(
        inst_i[2]), .C(n283), .ZN(n322) );
  OAI221V2_8TH40 U156 ( .A1(n276), .A2(n317), .B1(n278), .B2(n318), .C(n319), 
        .ZN(N1776) );
  AOI221V2_8TH40 U157 ( .A1(gpr2_data_i[19]), .A2(n281), .B1(n282), .B2(
        inst_i[3]), .C(n283), .ZN(n319) );
  OAI221V2_8TH40 U158 ( .A1(n276), .A2(n314), .B1(n278), .B2(n315), .C(n316), 
        .ZN(N1777) );
  AOI221V2_8TH40 U159 ( .A1(gpr2_data_i[20]), .A2(n281), .B1(n282), .B2(
        inst_i[4]), .C(n283), .ZN(n316) );
  OAI221V2_8TH40 U160 ( .A1(n276), .A2(n311), .B1(n278), .B2(n312), .C(n313), 
        .ZN(N1778) );
  AOI221V2_8TH40 U161 ( .A1(gpr2_data_i[21]), .A2(n281), .B1(n282), .B2(
        inst_i[5]), .C(n283), .ZN(n313) );
  OAI221V2_8TH40 U162 ( .A1(n276), .A2(n308), .B1(n278), .B2(n309), .C(n310), 
        .ZN(N1779) );
  AOI221V2_8TH40 U163 ( .A1(gpr2_data_i[22]), .A2(n281), .B1(n282), .B2(
        inst_i[6]), .C(n283), .ZN(n310) );
  OAI221V2_8TH40 U164 ( .A1(n276), .A2(n305), .B1(n278), .B2(n306), .C(n307), 
        .ZN(N1780) );
  AOI221V2_8TH40 U165 ( .A1(gpr2_data_i[23]), .A2(n281), .B1(n282), .B2(
        inst_i[7]), .C(n283), .ZN(n307) );
  OAI221V2_8TH40 U166 ( .A1(n276), .A2(n302), .B1(n278), .B2(n303), .C(n304), 
        .ZN(N1781) );
  AOI221V2_8TH40 U167 ( .A1(gpr2_data_i[24]), .A2(n281), .B1(n282), .B2(
        inst_i[8]), .C(n283), .ZN(n304) );
  OAI221V2_8TH40 U168 ( .A1(n276), .A2(n299), .B1(n278), .B2(n300), .C(n301), 
        .ZN(N1782) );
  AOI221V2_8TH40 U169 ( .A1(gpr2_data_i[25]), .A2(n281), .B1(n282), .B2(
        inst_i[9]), .C(n283), .ZN(n301) );
  OAI221V2_8TH40 U170 ( .A1(n276), .A2(n296), .B1(n278), .B2(n297), .C(n298), 
        .ZN(N1783) );
  AOI221V2_8TH40 U171 ( .A1(gpr2_data_i[26]), .A2(n281), .B1(n282), .B2(
        inst_i[10]), .C(n283), .ZN(n298) );
  OAI221V2_8TH40 U172 ( .A1(n276), .A2(n293), .B1(n278), .B2(n294), .C(n295), 
        .ZN(N1784) );
  AOI221V2_8TH40 U173 ( .A1(gpr2_data_i[27]), .A2(n281), .B1(n282), .B2(
        inst_i[11]), .C(n283), .ZN(n295) );
  OAI221V2_8TH40 U174 ( .A1(n276), .A2(n290), .B1(n278), .B2(n291), .C(n292), 
        .ZN(N1785) );
  AOI221V2_8TH40 U175 ( .A1(gpr2_data_i[28]), .A2(n281), .B1(n282), .B2(
        inst_i[12]), .C(n283), .ZN(n292) );
  OAI221V2_8TH40 U176 ( .A1(n276), .A2(n287), .B1(n278), .B2(n288), .C(n289), 
        .ZN(N1786) );
  AOI221V2_8TH40 U177 ( .A1(gpr2_data_i[29]), .A2(n281), .B1(n282), .B2(
        inst_i[13]), .C(n283), .ZN(n289) );
  OAI221V2_8TH40 U178 ( .A1(n276), .A2(n284), .B1(n278), .B2(n285), .C(n286), 
        .ZN(N1787) );
  AOI221V2_8TH40 U179 ( .A1(gpr2_data_i[30]), .A2(n281), .B1(n282), .B2(
        inst_i[14]), .C(n283), .ZN(n286) );
  OAI221V2_8TH40 U180 ( .A1(n276), .A2(n277), .B1(n278), .B2(n279), .C(n280), 
        .ZN(N1788) );
  AOI221V2_8TH40 U181 ( .A1(gpr2_data_i[31]), .A2(n281), .B1(n282), .B2(
        inst_i[15]), .C(n283), .ZN(n280) );
  I2NOR4V2_8TH40 U182 ( .A1(n462), .A2(n151), .B1(inst_i[20]), .B2(n463), .ZN(
        n100) );
  NAND4V2_8TH40 U183 ( .A1(n251), .A2(n252), .A3(n447), .A4(n158), .ZN(n125)
         );
  NAND4V2_8TH40 U184 ( .A1(n44), .A2(n42), .A3(n448), .A4(n449), .ZN(n447) );
  OAI22V2_8TH40 U185 ( .A1(n147), .A2(n148), .B1(n149), .B2(n150), .ZN(n114)
         );
  OAI211V2_8TH40 U186 ( .A1(n138), .A2(n139), .B(n140), .C(n141), .ZN(n130) );
  NAND4V2_8TH40 U187 ( .A1(n344), .A2(n158), .A3(n129), .A4(n507), .ZN(n244)
         );
  NAND4V2_8TH40 U188 ( .A1(df_exid_gpr_we), .A2(n483), .A3(n484), .A4(n485), 
        .ZN(n444) );
  NOR3V2_8TH40 U189 ( .A1(n486), .A2(n487), .A3(n488), .ZN(n485) );
  OAI211V2_8TH40 U190 ( .A1(n440), .A2(n404), .B(n441), .C(n442), .ZN(N1699)
         );
  AOI22V2_8TH40 U191 ( .A1(n399), .A2(df_exid_exe_result[0]), .B1(
        gpr1_data_i[0]), .B2(n401), .ZN(n442) );
  OAI211V2_8TH40 U192 ( .A1(n437), .A2(n404), .B(n438), .C(n439), .ZN(N1700)
         );
  AOI22V2_8TH40 U193 ( .A1(n399), .A2(df_exid_exe_result[1]), .B1(
        gpr1_data_i[1]), .B2(n401), .ZN(n439) );
  OAI211V2_8TH40 U194 ( .A1(n434), .A2(n404), .B(n435), .C(n436), .ZN(N1701)
         );
  AOI22V2_8TH40 U195 ( .A1(n399), .A2(df_exid_exe_result[2]), .B1(
        gpr1_data_i[2]), .B2(n401), .ZN(n436) );
  OAI211V2_8TH40 U196 ( .A1(n431), .A2(n404), .B(n432), .C(n433), .ZN(N1702)
         );
  AOI22V2_8TH40 U197 ( .A1(n399), .A2(df_exid_exe_result[3]), .B1(
        gpr1_data_i[3]), .B2(n401), .ZN(n433) );
  OAI211V2_8TH40 U198 ( .A1(n426), .A2(n404), .B(n427), .C(n428), .ZN(N1703)
         );
  AOI22V2_8TH40 U199 ( .A1(n399), .A2(df_exid_exe_result[4]), .B1(
        gpr1_data_i[4]), .B2(n401), .ZN(n428) );
  AOI21V2_8TH40 U200 ( .A1(n266), .A2(n267), .B(gpr1_data_o[31]), .ZN(n265) );
  NOR4V2_8TH40 U201 ( .A1(n268), .A2(n269), .A3(n270), .A4(n271), .ZN(n267) );
  NOR4V2_8TH40 U202 ( .A1(n272), .A2(n273), .A3(n274), .A4(n275), .ZN(n266) );
  NAND4V2_8TH40 U203 ( .A1(n393), .A2(df_exid_gpr_we), .A3(n394), .A4(n395), 
        .ZN(n384) );
  NOR3V2_8TH40 U204 ( .A1(n396), .A2(n397), .A3(n398), .ZN(n395) );
  AOI31V2_8TH40 U205 ( .A1(n84), .A2(n85), .A3(n86), .B(n87), .ZN(n83) );
  MOAI22V2_8TH40 U206 ( .A1(n171), .A2(n87), .B1(inst_i[17]), .B2(n100), .ZN(
        n168) );
  I2NOR3V2_8TH40 U207 ( .A1(n162), .A2(n85), .B(n172), .ZN(n171) );
  NAND4V2_8TH40 U208 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(n230)
         );
  NAND4V2_8TH40 U209 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(n229)
         );
  XOR2V0_8TH40 U210 ( .A1(df_exid_target_gpr[2]), .A2(gpr2_addr[2]), .Z(n397)
         );
  AOI31V2_8TH40 U211 ( .A1(n251), .A2(n252), .A3(n253), .B(rst), .ZN(n250) );
  AOI31V2_8TH40 U212 ( .A1(n126), .A2(n254), .A3(n239), .B(inst_i[5]), .ZN(
        n253) );
  AO222V2_8TH40 U213 ( .A1(gpr1_data_o[31]), .A2(n206), .B1(pc_plus4[31]), 
        .B2(n205), .C1(n4), .C2(n258), .Z(branch_target_addr[31]) );
  AO222V2_8TH40 U214 ( .A1(gpr1_data_o[30]), .A2(n206), .B1(pc_plus4[30]), 
        .B2(n205), .C1(n5), .C2(n258), .Z(branch_target_addr[30]) );
  AO222V2_8TH40 U215 ( .A1(gpr1_data_o[29]), .A2(n206), .B1(pc_plus4[29]), 
        .B2(n205), .C1(n6), .C2(n258), .Z(branch_target_addr[29]) );
  AO222V2_8TH40 U216 ( .A1(gpr1_data_o[28]), .A2(n206), .B1(pc_plus4[28]), 
        .B2(n205), .C1(n7), .C2(n258), .Z(branch_target_addr[28]) );
  AO222V2_8TH40 U217 ( .A1(gpr1_data_o[27]), .A2(n206), .B1(n205), .B2(
        inst_i[25]), .C1(n8), .C2(n258), .Z(branch_target_addr[27]) );
  AO222V2_8TH40 U218 ( .A1(gpr1_data_o[26]), .A2(n206), .B1(n205), .B2(
        inst_i[24]), .C1(n9), .C2(n258), .Z(branch_target_addr[26]) );
  AO222V2_8TH40 U219 ( .A1(gpr1_data_o[25]), .A2(n206), .B1(n205), .B2(
        inst_i[23]), .C1(n10), .C2(n258), .Z(branch_target_addr[25]) );
  AO222V2_8TH40 U220 ( .A1(gpr1_data_o[24]), .A2(n206), .B1(n205), .B2(
        inst_i[22]), .C1(n11), .C2(n258), .Z(branch_target_addr[24]) );
  AO222V2_8TH40 U221 ( .A1(gpr1_data_o[23]), .A2(n206), .B1(n205), .B2(
        inst_i[21]), .C1(n12), .C2(n258), .Z(branch_target_addr[23]) );
  AO222V2_8TH40 U222 ( .A1(n13), .A2(n258), .B1(gpr1_data_o[22]), .B2(n206), 
        .C1(gpr2_addr[4]), .C2(n259), .Z(branch_target_addr[22]) );
  AO222V2_8TH40 U223 ( .A1(n16), .A2(n258), .B1(gpr1_data_o[19]), .B2(n206), 
        .C1(gpr2_addr[1]), .C2(n259), .Z(branch_target_addr[19]) );
  AO222V2_8TH40 U224 ( .A1(n17), .A2(n258), .B1(gpr1_data_o[18]), .B2(n206), 
        .C1(gpr2_addr[0]), .C2(n259), .Z(branch_target_addr[18]) );
  AO222V2_8TH40 U225 ( .A1(gpr1_data_o[17]), .A2(n206), .B1(n205), .B2(
        inst_i[15]), .C1(n18), .C2(n258), .Z(branch_target_addr[17]) );
  AO222V2_8TH40 U226 ( .A1(gpr1_data_o[16]), .A2(n206), .B1(n205), .B2(
        inst_i[14]), .C1(n19), .C2(n258), .Z(branch_target_addr[16]) );
  AO222V2_8TH40 U227 ( .A1(gpr1_data_o[15]), .A2(n206), .B1(n205), .B2(
        inst_i[13]), .C1(n20), .C2(n258), .Z(branch_target_addr[15]) );
  AO222V2_8TH40 U228 ( .A1(gpr1_data_o[14]), .A2(n206), .B1(n205), .B2(
        inst_i[12]), .C1(n21), .C2(n258), .Z(branch_target_addr[14]) );
  AO222V2_8TH40 U229 ( .A1(gpr1_data_o[13]), .A2(n206), .B1(n205), .B2(
        inst_i[11]), .C1(n22), .C2(n258), .Z(branch_target_addr[13]) );
  AO222V2_8TH40 U230 ( .A1(gpr1_data_o[12]), .A2(n206), .B1(inst_i[10]), .B2(
        n205), .C1(n23), .C2(n258), .Z(branch_target_addr[12]) );
  AO222V2_8TH40 U231 ( .A1(gpr1_data_o[11]), .A2(n206), .B1(inst_i[9]), .B2(
        n205), .C1(n24), .C2(n258), .Z(branch_target_addr[11]) );
  AO222V2_8TH40 U232 ( .A1(gpr1_data_o[10]), .A2(n206), .B1(inst_i[8]), .B2(
        n205), .C1(n25), .C2(n258), .Z(branch_target_addr[10]) );
  AO222V2_8TH40 U233 ( .A1(gpr1_data_o[9]), .A2(n206), .B1(inst_i[7]), .B2(
        n205), .C1(n26), .C2(n258), .Z(branch_target_addr[9]) );
  AO222V2_8TH40 U234 ( .A1(gpr1_data_o[8]), .A2(n206), .B1(inst_i[6]), .B2(
        n205), .C1(n27), .C2(n258), .Z(branch_target_addr[8]) );
  AO222V2_8TH40 U235 ( .A1(gpr1_data_o[7]), .A2(n206), .B1(n205), .B2(
        inst_i[5]), .C1(n28), .C2(n258), .Z(branch_target_addr[7]) );
  AO222V2_8TH40 U236 ( .A1(gpr1_data_o[6]), .A2(n206), .B1(n205), .B2(
        inst_i[4]), .C1(n29), .C2(n258), .Z(branch_target_addr[6]) );
  AO222V2_8TH40 U237 ( .A1(gpr1_data_o[5]), .A2(n206), .B1(n205), .B2(
        inst_i[3]), .C1(n30), .C2(n258), .Z(branch_target_addr[5]) );
  AO222V2_8TH40 U238 ( .A1(gpr1_data_o[4]), .A2(n206), .B1(n205), .B2(
        inst_i[2]), .C1(n31), .C2(n258), .Z(branch_target_addr[4]) );
  AO222V2_8TH40 U239 ( .A1(gpr1_data_o[3]), .A2(n206), .B1(n205), .B2(
        inst_i[1]), .C1(n32), .C2(n258), .Z(branch_target_addr[3]) );
  AO222V2_8TH40 U240 ( .A1(gpr1_data_o[2]), .A2(n206), .B1(n205), .B2(
        inst_i[0]), .C1(n33), .C2(n258), .Z(branch_target_addr[2]) );
  AND4V2_8TH40 U241 ( .A1(n480), .A2(ex_inst_type[7]), .A3(ex_inst_type[6]), 
        .A4(ex_inst_type[5]), .Z(n392) );
  OAI32V2_8TH40 U242 ( .A1(n132), .A2(n133), .A3(n134), .B1(rst), .B2(n135), 
        .ZN(inst_type[1]) );
  NOR4V2_8TH40 U243 ( .A1(n136), .A2(n137), .A3(n114), .A4(n130), .ZN(n135) );
  OAI222V2_8TH40 U244 ( .A1(n152), .A2(n147), .B1(n153), .B2(n87), .C1(n154), 
        .C2(n155), .ZN(n136) );
  AOAI211V2_8TH40 U245 ( .A1(n218), .A2(n219), .B(rst), .C(n59), .ZN(gpr_we)
         );
  AOI211V2_8TH40 U246 ( .A1(n64), .A2(n222), .B(n80), .C(n170), .ZN(n219) );
  AOI21V2_8TH40 U247 ( .A1(n75), .A2(n76), .B(rst), .ZN(inst_type[4]) );
  INOR4V2_8TH40 U248 ( .A1(n61), .B1(n81), .B2(n82), .B3(n83), .ZN(n75) );
  AOI31V2_8TH40 U249 ( .A1(n165), .A2(n166), .A3(n167), .B(rst), .ZN(
        inst_type[0]) );
  NOR4V2_8TH40 U250 ( .A1(n168), .A2(n169), .A3(n78), .A4(n170), .ZN(n167) );
  AOI31V2_8TH40 U251 ( .A1(n115), .A2(n116), .A3(n117), .B(rst), .ZN(
        inst_type[2]) );
  AOI31V2_8TH40 U252 ( .A1(n97), .A2(n98), .A3(n99), .B(rst), .ZN(inst_type[3]) );
  AOAI211V2_8TH40 U253 ( .A1(n67), .A2(n68), .B(rst), .C(n69), .ZN(
        inst_type[5]) );
  I2NOR4V2_8TH40 U254 ( .A1(n246), .A2(n60), .B1(n247), .B2(n243), .ZN(
        except_type[9]) );
  AOAI211V2_8TH40 U255 ( .A1(n248), .A2(n249), .B(n87), .C(n250), .ZN(n247) );
  AOAI211V2_8TH40 U256 ( .A1(n202), .A2(n203), .B(rst), .C(n198), .ZN(
        inst_class[1]) );
  OAI211V2_8TH40 U257 ( .A1(rst), .A2(n197), .B(n69), .C(n198), .ZN(
        inst_class[2]) );
  AOI31V2_8TH40 U258 ( .A1(n60), .A2(n61), .A3(n62), .B(rst), .ZN(inst_type[6]) );
  AOI31V2_8TH40 U259 ( .A1(n208), .A2(n77), .A3(n209), .B(rst), .ZN(
        inst_class[0]) );
  OAI221V0_8TH40 U260 ( .A1(n1), .A2(n2), .B1(n3), .B2(n40), .C(n41), .ZN(
        target_gpr[4]) );
  OAI221V0_8TH40 U261 ( .A1(n1), .A2(n42), .B1(n3), .B2(n43), .C(n41), .ZN(
        target_gpr[3]) );
  OAI221V0_8TH40 U262 ( .A1(n1), .A2(n44), .B1(n3), .B2(n45), .C(n41), .ZN(
        target_gpr[2]) );
  OAI221V0_8TH40 U263 ( .A1(n1), .A2(n46), .B1(n3), .B2(n47), .C(n41), .ZN(
        target_gpr[1]) );
  OAI221V0_8TH40 U264 ( .A1(n1), .A2(n48), .B1(n3), .B2(n49), .C(n41), .ZN(
        target_gpr[0]) );
  OR2V0_8TH40 U265 ( .A1(n50), .A2(rst), .Z(n41) );
  I2NAND4V0_8TH40 U266 ( .A1(n53), .A2(n54), .B1(n55), .B2(n56), .ZN(n52) );
  AOI21V0_8TH40 U267 ( .A1(n57), .A2(n58), .B(rst), .ZN(stall_req) );
  INOR2V0_8TH40 U268 ( .A1(pc_plus8[2]), .B1(n59), .ZN(link_addr[2]) );
  INOR2V0_8TH40 U269 ( .A1(pc_plus8[1]), .B1(n59), .ZN(link_addr[1]) );
  INOR2V0_8TH40 U270 ( .A1(pc_plus8[0]), .B1(n59), .ZN(link_addr[0]) );
  AOI211V0_8TH40 U271 ( .A1(n63), .A2(n64), .B(n65), .C(n66), .ZN(n62) );
  AOI211V0_8TH40 U272 ( .A1(n64), .A2(n70), .B(n71), .C(n72), .ZN(n68) );
  NOR2V0P5_8TH40 U273 ( .A1(n73), .A2(n74), .ZN(n67) );
  INOR4V0_8TH40 U274 ( .A1(n77), .B1(n78), .B2(n79), .B3(n80), .ZN(n76) );
  NOR4V0P5_8TH40 U275 ( .A1(n88), .A2(n89), .A3(n90), .A4(n63), .ZN(n86) );
  AOI22V0_8TH40 U276 ( .A1(n91), .A2(inst_i[5]), .B1(n92), .B2(n93), .ZN(n84)
         );
  AOI21V0_8TH40 U277 ( .A1(n94), .A2(n95), .B(n72), .ZN(n61) );
  CLKNV1_8TH40 U278 ( .I(n96), .ZN(n72) );
  NOR4V0P5_8TH40 U279 ( .A1(n105), .A2(n106), .A3(n88), .A4(n107), .ZN(n103)
         );
  NOR4V0P5_8TH40 U280 ( .A1(n108), .A2(n109), .A3(n63), .A4(n110), .ZN(n102)
         );
  AOI21V0_8TH40 U281 ( .A1(n111), .A2(n112), .B(n74), .ZN(n98) );
  NOR2V0P5_8TH40 U282 ( .A1(n113), .A2(n114), .ZN(n97) );
  AOI22V0_8TH40 U283 ( .A1(n121), .A2(n81), .B1(n122), .B2(n123), .ZN(n118) );
  IAO21V0_8TH40 U284 ( .A1(n87), .A2(n124), .B(n113), .ZN(n116) );
  OAI211V0_8TH40 U285 ( .A1(n125), .A2(n126), .B(n96), .C(n127), .ZN(n113) );
  CLKNAND2V1_8TH40 U286 ( .A1(n128), .A2(n129), .ZN(n96) );
  NOR2V0P5_8TH40 U287 ( .A1(n130), .A2(n131), .ZN(n115) );
  AOI22V0_8TH40 U288 ( .A1(n142), .A2(n93), .B1(n95), .B2(n143), .ZN(n141) );
  AOI31V0_8TH40 U289 ( .A1(n144), .A2(inst_i[28]), .A3(n145), .B(n146), .ZN(
        n140) );
  NOR2V0P5_8TH40 U290 ( .A1(inst_i[20]), .A2(n151), .ZN(n149) );
  NOR3V0P5_8TH40 U291 ( .A1(n158), .A2(n133), .A3(n134), .ZN(n157) );
  OAI211V0_8TH40 U292 ( .A1(n159), .A2(n160), .B(n161), .C(n162), .ZN(n156) );
  CLKNV1_8TH40 U293 ( .I(n163), .ZN(n152) );
  AND2V0_8TH40 U294 ( .A1(n160), .A2(n164), .Z(n133) );
  OAI222V0_8TH40 U295 ( .A1(n173), .A2(n174), .B1(n164), .B2(n175), .C1(n176), 
        .C2(n177), .ZN(n172) );
  OAOI211V0_8TH40 U296 ( .A1(n180), .A2(n181), .B(n159), .C(n160), .ZN(n179)
         );
  AOI31V0_8TH40 U297 ( .A1(inst_i[5]), .A2(n182), .A3(n183), .B(n110), .ZN(
        n162) );
  AOI222V0_8TH40 U298 ( .A1(n184), .A2(n111), .B1(n143), .B2(n163), .C1(n81), 
        .C2(n122), .ZN(n166) );
  INAND2V0_8TH40 U299 ( .A1(n185), .B1(n186), .ZN(n163) );
  NOR2V0P5_8TH40 U300 ( .A1(n131), .A2(n137), .ZN(n165) );
  OAI21V0_8TH40 U301 ( .A1(n145), .A2(n143), .B(n81), .ZN(n189) );
  AOI31V0_8TH40 U302 ( .A1(n128), .A2(n182), .A3(n183), .B(n54), .ZN(n188) );
  AOI22V0_8TH40 U303 ( .A1(n190), .A2(n142), .B1(n121), .B2(n185), .ZN(n187)
         );
  IOA21V0_8TH40 U304 ( .A1(n191), .A2(n144), .B(n192), .ZN(n185) );
  OAI21V0_8TH40 U305 ( .A1(n193), .A2(n148), .B(n194), .ZN(n74) );
  AOI22V0_8TH40 U306 ( .A1(n123), .A2(n143), .B1(n95), .B2(n122), .ZN(n196) );
  CLKNV1_8TH40 U307 ( .I(n120), .ZN(n139) );
  CLKNV1_8TH40 U308 ( .I(inst_type[7]), .ZN(n69) );
  AOI21V0_8TH40 U309 ( .A1(n199), .A2(n200), .B(rst), .ZN(inst_type[7]) );
  IAO21V0_8TH40 U310 ( .A1(n87), .A2(n201), .B(n95), .ZN(n197) );
  AOI211V0_8TH40 U311 ( .A1(n51), .A2(n204), .B(n205), .C(n206), .ZN(n198) );
  CLKNV1_8TH40 U312 ( .I(n207), .ZN(n202) );
  AOI211V0_8TH40 U313 ( .A1(n210), .A2(n64), .B(n207), .C(n211), .ZN(n209) );
  OAI21V0_8TH40 U314 ( .A1(n106), .A2(n215), .B(n64), .ZN(n214) );
  NOR2V0P5_8TH40 U315 ( .A1(n216), .A2(n217), .ZN(n208) );
  AOI21V0_8TH40 U316 ( .A1(n169), .A2(inst_i[20]), .B(n79), .ZN(n50) );
  CLKNV1_8TH40 U317 ( .I(n178), .ZN(n221) );
  AND2V0_8TH40 U318 ( .A1(n142), .A2(n223), .Z(n170) );
  NOR2V0P5_8TH40 U319 ( .A1(n154), .A2(n164), .ZN(n142) );
  NOR2V0P5_8TH40 U320 ( .A1(n210), .A2(n226), .ZN(n225) );
  MUX2NV0_8TH40 U321 ( .I0(n227), .I1(n223), .S(n228), .ZN(n224) );
  NOR4V0P5_8TH40 U322 ( .A1(gpr2_data_o[23]), .A2(gpr2_data_o[22]), .A3(
        gpr2_data_o[21]), .A4(gpr2_data_o[20]), .ZN(n234) );
  NOR4V0P5_8TH40 U323 ( .A1(gpr2_data_o[1]), .A2(gpr2_data_o[19]), .A3(
        gpr2_data_o[18]), .A4(gpr2_data_o[17]), .ZN(n233) );
  NOR4V0P5_8TH40 U324 ( .A1(gpr2_data_o[16]), .A2(gpr2_data_o[15]), .A3(
        gpr2_data_o[14]), .A4(gpr2_data_o[13]), .ZN(n232) );
  NOR4V0P5_8TH40 U325 ( .A1(gpr2_data_o[12]), .A2(gpr2_data_o[11]), .A3(
        gpr2_data_o[10]), .A4(gpr2_data_o[0]), .ZN(n231) );
  NOR4V0P5_8TH40 U326 ( .A1(gpr2_data_o[9]), .A2(gpr2_data_o[8]), .A3(
        gpr2_data_o[7]), .A4(gpr2_data_o[6]), .ZN(n238) );
  NOR4V0P5_8TH40 U327 ( .A1(gpr2_data_o[5]), .A2(gpr2_data_o[4]), .A3(
        gpr2_data_o[3]), .A4(gpr2_data_o[31]), .ZN(n237) );
  NOR4V0P5_8TH40 U328 ( .A1(gpr2_data_o[30]), .A2(gpr2_data_o[2]), .A3(
        gpr2_data_o[29]), .A4(gpr2_data_o[28]), .ZN(n236) );
  NOR4V0P5_8TH40 U329 ( .A1(gpr2_data_o[27]), .A2(gpr2_data_o[26]), .A3(
        gpr2_data_o[25]), .A4(gpr2_data_o[24]), .ZN(n235) );
  AND2V0_8TH40 U330 ( .A1(n3), .A2(n203), .Z(n218) );
  CLKNAND2V1_8TH40 U331 ( .A1(n91), .A2(n128), .ZN(n77) );
  AOAI211V0_8TH40 U332 ( .A1(n241), .A2(n158), .B(n63), .C(n64), .ZN(n240) );
  INOR4V0_8TH40 U333 ( .A1(n242), .B1(n243), .B2(n73), .B3(n78), .ZN(n3) );
  NOR3V0P5_8TH40 U334 ( .A1(n212), .A2(n244), .A3(n245), .ZN(n78) );
  NOR2V0P5_8TH40 U335 ( .A1(rst), .A2(n194), .ZN(except_type[12]) );
  CLKNV1_8TH40 U336 ( .I(n91), .ZN(n254) );
  OAOI211V0_8TH40 U337 ( .A1(n181), .A2(inst_i[0]), .B(n134), .C(n160), .ZN(
        n91) );
  CLKNV1_8TH40 U338 ( .I(n226), .ZN(n249) );
  OA211V0_8TH40 U339 ( .A1(n212), .A2(n213), .B(n194), .C(n255), .Z(n60) );
  NAND4V0P5_8TH40 U340 ( .A1(n92), .A2(n93), .A3(inst_i[25]), .A4(n256), .ZN(
        n194) );
  NOR2V0P5_8TH40 U341 ( .A1(n126), .A2(n132), .ZN(except_type[8]) );
  INAND3V0_8TH40 U342 ( .A1(n177), .B1(n257), .B2(n180), .ZN(n126) );
  INOR2V0_8TH40 U343 ( .A1(curid_inst_delayslot_i), .B1(rst), .ZN(
        curid_inst_delayslot_o) );
  AO222V0_8TH40 U344 ( .A1(n14), .A2(n258), .B1(gpr1_data_o[21]), .B2(n206), 
        .C1(gpr2_addr[3]), .C2(n259), .Z(branch_target_addr[21]) );
  AO222V0_8TH40 U345 ( .A1(n15), .A2(n258), .B1(gpr1_data_o[20]), .B2(n206), 
        .C1(gpr2_addr[2]), .C2(n259), .Z(branch_target_addr[20]) );
  AO22V0_8TH40 U346 ( .A1(n206), .A2(gpr1_data_o[1]), .B1(n34), .B2(n258), .Z(
        branch_target_addr[1]) );
  AO22V0_8TH40 U347 ( .A1(n206), .A2(gpr1_data_o[0]), .B1(n35), .B2(n258), .Z(
        branch_target_addr[0]) );
  OR3V0_8TH40 U348 ( .A1(n205), .A2(n206), .A3(n258), .Z(branch_flag) );
  MUX2NV0_8TH40 U349 ( .I0(n145), .I1(n121), .S(n265), .ZN(n263) );
  OR4V0_8TH40 U350 ( .A1(gpr1_data_o[23]), .A2(gpr1_data_o[24]), .A3(
        gpr1_data_o[25]), .A4(gpr1_data_o[26]), .Z(n271) );
  OR4V0_8TH40 U351 ( .A1(gpr1_data_o[27]), .A2(gpr1_data_o[28]), .A3(
        gpr1_data_o[29]), .A4(gpr1_data_o[2]), .Z(n270) );
  OR4V0_8TH40 U352 ( .A1(gpr1_data_o[30]), .A2(gpr1_data_o[3]), .A3(
        gpr1_data_o[4]), .A4(gpr1_data_o[5]), .Z(n269) );
  OR4V0_8TH40 U353 ( .A1(gpr1_data_o[6]), .A2(gpr1_data_o[7]), .A3(
        gpr1_data_o[8]), .A4(gpr1_data_o[9]), .Z(n268) );
  OR3V0_8TH40 U354 ( .A1(gpr1_data_o[10]), .A2(gpr1_data_o[11]), .A3(
        gpr1_data_o[0]), .Z(n275) );
  OR4V0_8TH40 U355 ( .A1(gpr1_data_o[12]), .A2(gpr1_data_o[13]), .A3(
        gpr1_data_o[14]), .A4(gpr1_data_o[15]), .Z(n274) );
  OR4V0_8TH40 U356 ( .A1(gpr1_data_o[16]), .A2(gpr1_data_o[17]), .A3(
        gpr1_data_o[18]), .A4(gpr1_data_o[19]), .Z(n273) );
  OR4V0_8TH40 U357 ( .A1(gpr1_data_o[1]), .A2(gpr1_data_o[20]), .A3(
        gpr1_data_o[21]), .A4(gpr1_data_o[22]), .Z(n272) );
  MUX2NV0_8TH40 U358 ( .I0(n143), .I1(n122), .S(N812), .ZN(n262) );
  CLKXOR2V2_8TH40 U359 ( .A1(inst_i[16]), .A2(gpr1_data_o[31]), .Z(n260) );
  I2NOR3V1_8TH40 U360 ( .A1(n64), .A2(n108), .B(rst), .ZN(n206) );
  CLKNV1_8TH40 U361 ( .I(n87), .ZN(n64) );
  NOR2V0P5_8TH40 U362 ( .A1(rst), .A2(n255), .ZN(n205) );
  CLKNV1_8TH40 U363 ( .I(df_exid_exe_result[31]), .ZN(n279) );
  CLKNV1_8TH40 U364 ( .I(df_memid_exe_result[31]), .ZN(n277) );
  CLKNV1_8TH40 U365 ( .I(df_exid_exe_result[30]), .ZN(n285) );
  CLKNV1_8TH40 U366 ( .I(df_memid_exe_result[30]), .ZN(n284) );
  CLKNV1_8TH40 U367 ( .I(df_exid_exe_result[29]), .ZN(n288) );
  CLKNV1_8TH40 U368 ( .I(df_memid_exe_result[29]), .ZN(n287) );
  CLKNV1_8TH40 U369 ( .I(df_exid_exe_result[28]), .ZN(n291) );
  CLKNV1_8TH40 U370 ( .I(df_memid_exe_result[28]), .ZN(n290) );
  CLKNV1_8TH40 U371 ( .I(df_exid_exe_result[27]), .ZN(n294) );
  CLKNV1_8TH40 U372 ( .I(df_memid_exe_result[27]), .ZN(n293) );
  CLKNV1_8TH40 U373 ( .I(df_exid_exe_result[26]), .ZN(n297) );
  CLKNV1_8TH40 U374 ( .I(df_memid_exe_result[26]), .ZN(n296) );
  CLKNV1_8TH40 U375 ( .I(df_exid_exe_result[25]), .ZN(n300) );
  CLKNV1_8TH40 U376 ( .I(df_memid_exe_result[25]), .ZN(n299) );
  CLKNV1_8TH40 U377 ( .I(df_exid_exe_result[24]), .ZN(n303) );
  CLKNV1_8TH40 U378 ( .I(df_memid_exe_result[24]), .ZN(n302) );
  CLKNV1_8TH40 U379 ( .I(df_exid_exe_result[23]), .ZN(n306) );
  CLKNV1_8TH40 U380 ( .I(df_memid_exe_result[23]), .ZN(n305) );
  CLKNV1_8TH40 U381 ( .I(df_exid_exe_result[22]), .ZN(n309) );
  CLKNV1_8TH40 U382 ( .I(df_memid_exe_result[22]), .ZN(n308) );
  CLKNV1_8TH40 U383 ( .I(df_exid_exe_result[21]), .ZN(n312) );
  CLKNV1_8TH40 U384 ( .I(df_memid_exe_result[21]), .ZN(n311) );
  CLKNV1_8TH40 U385 ( .I(df_exid_exe_result[20]), .ZN(n315) );
  CLKNV1_8TH40 U386 ( .I(df_memid_exe_result[20]), .ZN(n314) );
  CLKNV1_8TH40 U387 ( .I(df_exid_exe_result[19]), .ZN(n318) );
  CLKNV1_8TH40 U388 ( .I(df_memid_exe_result[19]), .ZN(n317) );
  CLKNV1_8TH40 U389 ( .I(df_exid_exe_result[18]), .ZN(n321) );
  CLKNV1_8TH40 U390 ( .I(df_memid_exe_result[18]), .ZN(n320) );
  CLKNV1_8TH40 U391 ( .I(df_exid_exe_result[17]), .ZN(n324) );
  CLKNV1_8TH40 U392 ( .I(df_memid_exe_result[17]), .ZN(n323) );
  I2NOR4V0_8TH40 U393 ( .A1(n329), .A2(n330), .B1(n2), .B2(rst), .ZN(n283) );
  NOR3V0P5_8TH40 U394 ( .A1(n331), .A2(rst), .A3(n195), .ZN(n282) );
  CLKNV1_8TH40 U395 ( .I(df_exid_exe_result[16]), .ZN(n327) );
  CLKNV1_8TH40 U396 ( .I(df_memid_exe_result[16]), .ZN(n326) );
  CLKNV1_8TH40 U397 ( .I(n332), .ZN(n276) );
  CLKNV1_8TH40 U398 ( .I(df_exid_exe_result[15]), .ZN(n334) );
  CLKNV1_8TH40 U399 ( .I(df_exid_exe_result[14]), .ZN(n336) );
  CLKNV1_8TH40 U400 ( .I(df_exid_exe_result[13]), .ZN(n338) );
  CLKNV1_8TH40 U401 ( .I(df_exid_exe_result[12]), .ZN(n340) );
  CLKNV1_8TH40 U402 ( .I(df_exid_exe_result[11]), .ZN(n342) );
  CLKNV1_8TH40 U403 ( .I(df_exid_exe_result[10]), .ZN(n345) );
  CLKNV1_8TH40 U404 ( .I(df_exid_exe_result[9]), .ZN(n348) );
  CLKNV1_8TH40 U405 ( .I(df_exid_exe_result[8]), .ZN(n351) );
  CLKNV1_8TH40 U406 ( .I(df_exid_exe_result[7]), .ZN(n354) );
  CLKNV1_8TH40 U407 ( .I(df_exid_exe_result[6]), .ZN(n357) );
  CLKNV1_8TH40 U408 ( .I(df_exid_exe_result[5]), .ZN(n359) );
  CLKNV1_8TH40 U409 ( .I(df_exid_exe_result[4]), .ZN(n362) );
  CLKNV1_8TH40 U410 ( .I(df_exid_exe_result[3]), .ZN(n365) );
  CLKNV1_8TH40 U411 ( .I(df_exid_exe_result[2]), .ZN(n368) );
  CLKNV1_8TH40 U412 ( .I(df_exid_exe_result[1]), .ZN(n371) );
  NOR2V0P5_8TH40 U413 ( .A1(n375), .A2(n331), .ZN(n332) );
  I2NOR3V1_8TH40 U414 ( .A1(gpr2_re), .A2(n375), .B(n331), .ZN(n281) );
  CLKXOR2V2_8TH40 U415 ( .A1(df_memid_target_gpr[4]), .A2(gpr2_addr[4]), .Z(
        n382) );
  CLKXOR2V2_8TH40 U416 ( .A1(df_memid_target_gpr[0]), .A2(n49), .Z(n378) );
  CLKXOR2V2_8TH40 U417 ( .A1(df_memid_target_gpr[2]), .A2(n45), .Z(n377) );
  CLKXOR2V2_8TH40 U418 ( .A1(df_memid_target_gpr[1]), .A2(n47), .Z(n376) );
  CLKNV1_8TH40 U419 ( .I(df_exid_exe_result[0]), .ZN(n373) );
  CLKNAND2V1_8TH40 U420 ( .A1(n383), .A2(n329), .ZN(n333) );
  CLKNV1_8TH40 U421 ( .I(n331), .ZN(n329) );
  NAND3V0P5_8TH40 U422 ( .A1(n278), .A2(n51), .A3(n331), .ZN(N1756) );
  OAI21V0_8TH40 U423 ( .A1(n384), .A2(n380), .B(n58), .ZN(n331) );
  NAND3V0P5_8TH40 U424 ( .A1(n385), .A2(n58), .A3(gpr2_re), .ZN(n278) );
  CLKNV1_8TH40 U425 ( .I(n380), .ZN(gpr2_re) );
  INOR4V0_8TH40 U426 ( .A1(n161), .B1(n226), .B2(n105), .B3(n70), .ZN(n389) );
  NOR4V0P5_8TH40 U427 ( .A1(n177), .A2(n370), .A3(n173), .A4(n367), .ZN(n226)
         );
  OAI21V0_8TH40 U428 ( .A1(n264), .A2(n391), .B(n104), .ZN(n390) );
  CLKNAND2V1_8TH40 U429 ( .A1(n82), .A2(inst_i[29]), .ZN(n104) );
  CLKNAND2V1_8TH40 U430 ( .A1(n392), .A2(n385), .ZN(n58) );
  CLKNV1_8TH40 U431 ( .I(n384), .ZN(n385) );
  CLKXOR2V2_8TH40 U432 ( .A1(df_exid_target_gpr[1]), .A2(gpr2_addr[1]), .Z(
        n398) );
  CLKXOR2V2_8TH40 U433 ( .A1(df_exid_target_gpr[0]), .A2(gpr2_addr[0]), .Z(
        n396) );
  CLKXOR2V2_8TH40 U434 ( .A1(df_exid_target_gpr[3]), .A2(n43), .Z(n394) );
  CLKXOR2V2_8TH40 U435 ( .A1(df_exid_target_gpr[4]), .A2(n40), .Z(n393) );
  CLKNV1_8TH40 U436 ( .I(df_memid_exe_result[15]), .ZN(n403) );
  CLKNV1_8TH40 U437 ( .I(inst_i[15]), .ZN(n2) );
  CLKNV1_8TH40 U438 ( .I(df_memid_exe_result[14]), .ZN(n406) );
  CLKNV1_8TH40 U439 ( .I(df_memid_exe_result[13]), .ZN(n408) );
  CLKNV1_8TH40 U440 ( .I(df_memid_exe_result[12]), .ZN(n410) );
  CLKNV1_8TH40 U441 ( .I(inst_i[12]), .ZN(n46) );
  CLKNV1_8TH40 U442 ( .I(df_memid_exe_result[11]), .ZN(n412) );
  CLKNV1_8TH40 U443 ( .I(inst_i[11]), .ZN(n48) );
  CLKNV1_8TH40 U444 ( .I(df_memid_exe_result[10]), .ZN(n414) );
  CLKNV1_8TH40 U445 ( .I(df_memid_exe_result[9]), .ZN(n416) );
  CLKNV1_8TH40 U446 ( .I(inst_i[9]), .ZN(n347) );
  CLKNV1_8TH40 U447 ( .I(df_memid_exe_result[8]), .ZN(n418) );
  CLKNV1_8TH40 U448 ( .I(inst_i[8]), .ZN(n350) );
  CLKNV1_8TH40 U449 ( .I(df_memid_exe_result[7]), .ZN(n420) );
  CLKNV1_8TH40 U450 ( .I(inst_i[7]), .ZN(n353) );
  CLKNV1_8TH40 U451 ( .I(df_memid_exe_result[6]), .ZN(n422) );
  CLKNV1_8TH40 U452 ( .I(inst_i[6]), .ZN(n356) );
  CLKNV1_8TH40 U453 ( .I(df_memid_exe_result[5]), .ZN(n424) );
  AOI22V0_8TH40 U454 ( .A1(n429), .A2(inst_i[4]), .B1(n430), .B2(inst_i[10]), 
        .ZN(n427) );
  CLKNV1_8TH40 U455 ( .I(df_memid_exe_result[4]), .ZN(n426) );
  AOI22V0_8TH40 U456 ( .A1(n429), .A2(inst_i[3]), .B1(n430), .B2(inst_i[9]), 
        .ZN(n432) );
  CLKNV1_8TH40 U457 ( .I(df_memid_exe_result[3]), .ZN(n431) );
  AOI22V0_8TH40 U458 ( .A1(n429), .A2(inst_i[2]), .B1(n430), .B2(inst_i[8]), 
        .ZN(n435) );
  CLKNV1_8TH40 U459 ( .I(df_memid_exe_result[2]), .ZN(n434) );
  AOI22V0_8TH40 U460 ( .A1(n429), .A2(inst_i[1]), .B1(n430), .B2(inst_i[7]), 
        .ZN(n438) );
  CLKNV1_8TH40 U461 ( .I(df_memid_exe_result[1]), .ZN(n437) );
  I2NOR3V1_8TH40 U462 ( .A1(n443), .A2(n444), .B(n445), .ZN(n401) );
  AOI22V0_8TH40 U463 ( .A1(n429), .A2(inst_i[0]), .B1(n430), .B2(inst_i[6]), 
        .ZN(n441) );
  NOR3V0P5_8TH40 U464 ( .A1(n446), .A2(n239), .A3(n132), .ZN(n430) );
  CLKNAND2V1_8TH40 U465 ( .A1(n128), .A2(n51), .ZN(n132) );
  CLKNV1_8TH40 U466 ( .I(n125), .ZN(n128) );
  NOR4V0P5_8TH40 U467 ( .A1(inst_i[12]), .A2(inst_i[11]), .A3(n450), .A4(n244), 
        .ZN(n449) );
  NOR3V0P5_8TH40 U468 ( .A1(inst_i[15]), .A2(inst_i[20]), .A3(inst_i[16]), 
        .ZN(n448) );
  CLKNV1_8TH40 U469 ( .I(inst_i[14]), .ZN(n42) );
  CLKNV1_8TH40 U470 ( .I(inst_i[13]), .ZN(n44) );
  CLKNV1_8TH40 U471 ( .I(n245), .ZN(n252) );
  CLKNV1_8TH40 U472 ( .I(n402), .ZN(n429) );
  NAND3V0P5_8TH40 U473 ( .A1(n57), .A2(n445), .A3(n383), .ZN(n402) );
  OA31V0_8TH40 U474 ( .A1(n330), .A2(n217), .A3(n451), .B(n51), .Z(n383) );
  CLKNAND2V1_8TH40 U475 ( .A1(n452), .A2(n148), .ZN(n330) );
  CLKNV1_8TH40 U476 ( .I(n400), .ZN(n404) );
  NOR2V0P5_8TH40 U477 ( .A1(n443), .A2(n453), .ZN(n400) );
  CLKXOR2V2_8TH40 U478 ( .A1(gpr1_addr[4]), .A2(df_memid_target_gpr[4]), .Z(
        n459) );
  CLKXOR2V2_8TH40 U479 ( .A1(gpr1_addr[1]), .A2(df_memid_target_gpr[1]), .Z(
        n458) );
  CLKXOR2V2_8TH40 U480 ( .A1(gpr1_addr[0]), .A2(df_memid_target_gpr[0]), .Z(
        n457) );
  CLKNV1_8TH40 U481 ( .I(n460), .ZN(gpr1_addr[0]) );
  CLKXOR2V2_8TH40 U482 ( .A1(gpr1_addr[3]), .A2(df_memid_target_gpr[3]), .Z(
        n456) );
  XNOR2V0_8TH40 U483 ( .A1(df_memid_target_gpr[2]), .A2(gpr1_addr[2]), .ZN(
        n454) );
  CLKNV1_8TH40 U484 ( .I(n445), .ZN(gpr1_re) );
  CLKNV1_8TH40 U485 ( .I(n148), .ZN(n95) );
  OAI21V0_8TH40 U486 ( .A1(n248), .A2(n87), .B(n246), .ZN(n461) );
  I2NOR4V0_8TH40 U487 ( .A1(n200), .A2(n199), .B1(n65), .B2(n73), .ZN(n246) );
  OAI211V0_8TH40 U488 ( .A1(n147), .A2(n148), .B(n119), .C(n195), .ZN(n73) );
  INAND2V0_8TH40 U489 ( .A1(n204), .B1(n452), .ZN(n65) );
  NOR2V0P5_8TH40 U490 ( .A1(n120), .A2(n100), .ZN(n452) );
  CLKNV1_8TH40 U491 ( .I(inst_i[16]), .ZN(n151) );
  NOR2V0P5_8TH40 U492 ( .A1(n464), .A2(n465), .ZN(n462) );
  NOR4V0P5_8TH40 U493 ( .A1(n464), .A2(n463), .A3(inst_i[18]), .A4(inst_i[20]), 
        .ZN(n120) );
  CLKNAND2V1_8TH40 U494 ( .A1(n264), .A2(n150), .ZN(n204) );
  CLKNV1_8TH40 U495 ( .I(n169), .ZN(n150) );
  NOR2V0P5_8TH40 U496 ( .A1(n463), .A2(n450), .ZN(n169) );
  NAND3V0P5_8TH40 U497 ( .A1(n465), .A2(n464), .A3(n138), .ZN(n450) );
  CLKNV1_8TH40 U498 ( .I(inst_i[17]), .ZN(n138) );
  CLKNV1_8TH40 U499 ( .I(inst_i[19]), .ZN(n464) );
  CLKNV1_8TH40 U500 ( .I(inst_i[18]), .ZN(n465) );
  CLKNV1_8TH40 U501 ( .I(n66), .ZN(n199) );
  NOR2V0P5_8TH40 U502 ( .A1(n211), .A2(n80), .ZN(n200) );
  AND2V0_8TH40 U503 ( .A1(n466), .A2(n111), .Z(n80) );
  CLKNV1_8TH40 U504 ( .I(n184), .ZN(n468) );
  AOA211V0_8TH40 U505 ( .A1(n93), .A2(n182), .B(n112), .C(n111), .Z(n211) );
  CLKNV1_8TH40 U506 ( .I(n154), .ZN(n111) );
  NAND3V0P5_8TH40 U507 ( .A1(inst_i[28]), .A2(inst_i[29]), .A3(n469), .ZN(n154) );
  OAI31V0_8TH40 U508 ( .A1(n223), .A2(n178), .A3(n190), .B(n182), .ZN(n470) );
  NOR2V0P5_8TH40 U509 ( .A1(n173), .A2(n471), .ZN(n190) );
  CLKNAND2V1_8TH40 U510 ( .A1(n251), .A2(n245), .ZN(n87) );
  CLKNAND2V1_8TH40 U511 ( .A1(n472), .A2(n473), .ZN(n245) );
  NOR4V0P5_8TH40 U512 ( .A1(n63), .A2(n90), .A3(n89), .A4(n210), .ZN(n124) );
  CLKNAND2V1_8TH40 U513 ( .A1(n182), .A2(n257), .ZN(n476) );
  NOR3V0P5_8TH40 U514 ( .A1(n467), .A2(n471), .A3(n160), .ZN(n89) );
  NOR4V0P5_8TH40 U515 ( .A1(n160), .A2(n467), .A3(n370), .A4(n367), .ZN(n90)
         );
  CLKNAND2V1_8TH40 U516 ( .A1(inst_i[5]), .A2(n180), .ZN(n467) );
  CLKNV1_8TH40 U517 ( .I(n155), .ZN(n63) );
  NAND4V0P5_8TH40 U518 ( .A1(n257), .A2(n182), .A3(n180), .A4(n158), .ZN(n155)
         );
  CLKNV1_8TH40 U519 ( .I(n471), .ZN(n257) );
  CLKNAND2V1_8TH40 U520 ( .A1(inst_i[2]), .A2(n370), .ZN(n471) );
  INOR4V0_8TH40 U521 ( .A1(n477), .B1(n184), .B2(n110), .B3(n109), .ZN(n201)
         );
  NOR3V0P5_8TH40 U522 ( .A1(n177), .A2(n134), .A3(n158), .ZN(n109) );
  NOR3V0P5_8TH40 U523 ( .A1(n159), .A2(n177), .A3(n158), .ZN(n110) );
  NOR3V0P5_8TH40 U524 ( .A1(n164), .A2(n181), .A3(n175), .ZN(n184) );
  CLKNAND2V1_8TH40 U525 ( .A1(inst_i[5]), .A2(inst_i[0]), .ZN(n175) );
  INAND2V0_8TH40 U526 ( .A1(n239), .B1(inst_i[5]), .ZN(n477) );
  CLKNV1_8TH40 U527 ( .I(n134), .ZN(n478) );
  CLKNV1_8TH40 U528 ( .I(n159), .ZN(n183) );
  AO31V0_8TH40 U529 ( .A1(n159), .A2(n181), .A3(n134), .B(n158), .Z(n475) );
  NOR3V0P5_8TH40 U530 ( .A1(n108), .A2(n105), .A3(n215), .ZN(n474) );
  NOR2V0P5_8TH40 U531 ( .A1(n160), .A2(n176), .ZN(n215) );
  NOR2V0P5_8TH40 U532 ( .A1(n178), .A2(n227), .ZN(n176) );
  CLKNAND2V1_8TH40 U533 ( .A1(inst_i[4]), .A2(n364), .ZN(n160) );
  AND2V0_8TH40 U534 ( .A1(n479), .A2(n92), .Z(n105) );
  INOR2V0_8TH40 U535 ( .A1(n479), .B1(n177), .ZN(n108) );
  OR2V0_8TH40 U536 ( .A1(n93), .A2(n178), .Z(n479) );
  NOR2V0P5_8TH40 U537 ( .A1(n173), .A2(n181), .ZN(n178) );
  CLKNAND2V1_8TH40 U538 ( .A1(inst_i[0]), .A2(n158), .ZN(n173) );
  NOR3V0P5_8TH40 U539 ( .A1(inst_i[0]), .A2(inst_i[5]), .A3(n181), .ZN(n93) );
  NOR4V0P5_8TH40 U540 ( .A1(n241), .A2(n107), .A3(n88), .A4(n106), .ZN(n161)
         );
  IAO21V0_8TH40 U541 ( .A1(n227), .A2(n223), .B(n177), .ZN(n106) );
  CLKNAND2V1_8TH40 U542 ( .A1(inst_i[3]), .A2(n361), .ZN(n177) );
  AND2V0_8TH40 U543 ( .A1(n223), .A2(n92), .Z(n88) );
  NOR2V0P5_8TH40 U544 ( .A1(n134), .A2(inst_i[5]), .ZN(n223) );
  NAND3V0P5_8TH40 U545 ( .A1(n180), .A2(n367), .A3(inst_i[1]), .ZN(n134) );
  CLKNV1_8TH40 U546 ( .I(inst_i[0]), .ZN(n180) );
  AND2V0_8TH40 U547 ( .A1(n227), .A2(n92), .Z(n107) );
  NOR2V0P5_8TH40 U548 ( .A1(n361), .A2(n364), .ZN(n92) );
  NOR2V0P5_8TH40 U549 ( .A1(n159), .A2(inst_i[5]), .ZN(n227) );
  NAND3V0P5_8TH40 U550 ( .A1(inst_i[0]), .A2(n367), .A3(inst_i[1]), .ZN(n159)
         );
  CLKNV1_8TH40 U551 ( .I(n174), .ZN(n241) );
  NAND3V0P5_8TH40 U552 ( .A1(inst_i[2]), .A2(n182), .A3(inst_i[1]), .ZN(n174)
         );
  CLKNV1_8TH40 U553 ( .I(n164), .ZN(n182) );
  CLKNV1_8TH40 U554 ( .I(df_memid_exe_result[0]), .ZN(n440) );
  CLKNAND2V1_8TH40 U555 ( .A1(n446), .A2(n51), .ZN(N1698) );
  CLKNV1_8TH40 U556 ( .I(n57), .ZN(n446) );
  CLKNAND2V1_8TH40 U557 ( .A1(n453), .A2(n392), .ZN(n57) );
  OR3V0_8TH40 U558 ( .A1(ex_inst_type[1]), .A2(ex_inst_type[2]), .A3(
        ex_inst_type[0]), .Z(n482) );
  AO31V0_8TH40 U559 ( .A1(ex_inst_type[1]), .A2(ex_inst_type[0]), .A3(
        ex_inst_type[2]), .B(ex_inst_type[3]), .Z(n481) );
  CLKNV1_8TH40 U560 ( .I(n444), .ZN(n453) );
  CLKXOR2V2_8TH40 U561 ( .A1(gpr1_addr[4]), .A2(df_exid_target_gpr[4]), .Z(
        n488) );
  AO22V0_8TH40 U562 ( .A1(n489), .A2(inst_i[25]), .B1(gpr2_addr[4]), .B2(n71), 
        .Z(gpr1_addr[4]) );
  CLKNV1_8TH40 U563 ( .I(n40), .ZN(gpr2_addr[4]) );
  CLKNAND2V1_8TH40 U564 ( .A1(inst_i[20]), .A2(n51), .ZN(n40) );
  CLKXOR2V2_8TH40 U565 ( .A1(gpr1_addr[3]), .A2(df_exid_target_gpr[3]), .Z(
        n487) );
  CLKXOR2V2_8TH40 U566 ( .A1(gpr1_addr[1]), .A2(df_exid_target_gpr[1]), .Z(
        n486) );
  AO22V0_8TH40 U567 ( .A1(n489), .A2(inst_i[22]), .B1(gpr2_addr[1]), .B2(n71), 
        .Z(gpr1_addr[1]) );
  CLKNV1_8TH40 U568 ( .I(n47), .ZN(gpr2_addr[1]) );
  CLKNAND2V1_8TH40 U569 ( .A1(inst_i[17]), .A2(n51), .ZN(n47) );
  XNOR2V0_8TH40 U570 ( .A1(df_exid_target_gpr[2]), .A2(gpr1_addr[2]), .ZN(n484) );
  CLKNAND2V1_8TH40 U571 ( .A1(inst_i[18]), .A2(n51), .ZN(n45) );
  CLKXOR2V2_8TH40 U572 ( .A1(df_exid_target_gpr[0]), .A2(n460), .Z(n483) );
  AOI22V0_8TH40 U573 ( .A1(n489), .A2(inst_i[21]), .B1(gpr2_addr[0]), .B2(n71), 
        .ZN(n460) );
  INOR2V0_8TH40 U574 ( .A1(n53), .B1(n213), .ZN(n71) );
  NOR2V0P5_8TH40 U575 ( .A1(n473), .A2(n212), .ZN(n53) );
  CLKNV1_8TH40 U576 ( .I(inst_i[23]), .ZN(n473) );
  CLKNV1_8TH40 U577 ( .I(n49), .ZN(gpr2_addr[0]) );
  CLKNAND2V1_8TH40 U578 ( .A1(inst_i[16]), .A2(n51), .ZN(n49) );
  CLKNV1_8TH40 U579 ( .I(n490), .ZN(n489) );
  NOR3V0P5_8TH40 U580 ( .A1(n66), .A2(n243), .A3(n259), .ZN(n492) );
  CLKNV1_8TH40 U581 ( .I(n255), .ZN(n259) );
  NOR2V0P5_8TH40 U582 ( .A1(n54), .A2(n79), .ZN(n255) );
  AND2V0_8TH40 U583 ( .A1(n493), .A2(n121), .Z(n79) );
  CLKNV1_8TH40 U584 ( .I(n193), .ZN(n121) );
  CLKNV1_8TH40 U585 ( .I(n127), .ZN(n54) );
  CLKNAND2V1_8TH40 U586 ( .A1(n145), .A2(n493), .ZN(n127) );
  INAND2V0_8TH40 U587 ( .A1(n451), .B1(n148), .ZN(n243) );
  NAND3V0P5_8TH40 U588 ( .A1(n494), .A2(n191), .A3(inst_i[29]), .ZN(n148) );
  NOR4V0P5_8TH40 U589 ( .A1(n495), .A2(n496), .A3(n497), .A4(inst_i[28]), .ZN(
        n451) );
  CLKNAND2V1_8TH40 U590 ( .A1(n242), .A2(n56), .ZN(n66) );
  OAI21V0_8TH40 U591 ( .A1(n145), .A2(n191), .B(n144), .ZN(n56) );
  NOR3V0P5_8TH40 U592 ( .A1(n498), .A2(inst_i[30]), .A3(n499), .ZN(n144) );
  CLKNV1_8TH40 U593 ( .I(n147), .ZN(n145) );
  NOR4V0P5_8TH40 U594 ( .A1(n496), .A2(n501), .A3(n499), .A4(inst_i[28]), .ZN(
        n82) );
  AOI21V0_8TH40 U595 ( .A1(n123), .A2(n94), .B(n387), .ZN(n500) );
  IOAI21V1_8TH40 U596 ( .B1(n147), .B2(n192), .A(n146), .ZN(n387) );
  NOR4V0P5_8TH40 U597 ( .A1(n495), .A2(n191), .A3(inst_i[26]), .A4(inst_i[30]), 
        .ZN(n146) );
  CLKNV1_8TH40 U598 ( .I(n391), .ZN(n94) );
  NOR4V0P5_8TH40 U599 ( .A1(n191), .A2(n499), .A3(inst_i[29]), .A4(inst_i[30]), 
        .ZN(n123) );
  NAND3V0P5_8TH40 U600 ( .A1(n502), .A2(n496), .A3(inst_i[31]), .ZN(n192) );
  CLKNV1_8TH40 U601 ( .I(n264), .ZN(n81) );
  NAND3V0P5_8TH40 U602 ( .A1(n494), .A2(n498), .A3(inst_i[28]), .ZN(n264) );
  INOR2V0_8TH40 U603 ( .A1(n493), .B1(n501), .ZN(n251) );
  AOI22V0_8TH40 U604 ( .A1(inst_i[26]), .A2(n495), .B1(inst_i[29]), .B2(n499), 
        .ZN(n506) );
  NAND3V0P5_8TH40 U605 ( .A1(inst_i[27]), .A2(n498), .A3(inst_i[31]), .ZN(n495) );
  AOI211V0_8TH40 U606 ( .A1(n498), .A2(n193), .B(n191), .C(n499), .ZN(n504) );
  CLKNV1_8TH40 U607 ( .I(inst_i[31]), .ZN(n499) );
  CLKNV1_8TH40 U608 ( .I(inst_i[28]), .ZN(n191) );
  CLKNV1_8TH40 U609 ( .I(inst_i[29]), .ZN(n498) );
  INAND2V0_8TH40 U610 ( .A1(n244), .B1(n472), .ZN(n213) );
  NOR4V0P5_8TH40 U611 ( .A1(inst_i[21]), .A2(inst_i[22]), .A3(inst_i[24]), 
        .A4(inst_i[25]), .ZN(n472) );
  NOR4V0P5_8TH40 U612 ( .A1(inst_i[9]), .A2(inst_i[8]), .A3(inst_i[7]), .A4(
        inst_i[6]), .ZN(n507) );
  NOR3V0P5_8TH40 U613 ( .A1(n181), .A2(inst_i[0]), .A3(n164), .ZN(n129) );
  CLKNAND2V1_8TH40 U614 ( .A1(n361), .A2(n364), .ZN(n164) );
  CLKNV1_8TH40 U615 ( .I(inst_i[3]), .ZN(n364) );
  CLKNV1_8TH40 U616 ( .I(inst_i[4]), .ZN(n361) );
  CLKNAND2V1_8TH40 U617 ( .A1(n367), .A2(n370), .ZN(n181) );
  CLKNV1_8TH40 U618 ( .I(inst_i[1]), .ZN(n370) );
  CLKNV1_8TH40 U619 ( .I(inst_i[2]), .ZN(n367) );
  CLKNV1_8TH40 U620 ( .I(inst_i[5]), .ZN(n158) );
  CLKNV1_8TH40 U621 ( .I(inst_i[10]), .ZN(n344) );
  CLKNV1_8TH40 U622 ( .I(n212), .ZN(n256) );
  CLKNAND2V1_8TH40 U623 ( .A1(n469), .A2(n502), .ZN(n212) );
  NOR3V0P5_8TH40 U624 ( .A1(n501), .A2(inst_i[31]), .A3(n496), .ZN(n469) );
  CLKNV1_8TH40 U625 ( .I(inst_i[30]), .ZN(n496) );
  CLKNV1_8TH40 U626 ( .I(n122), .ZN(n501) );
  CLKNAND2V1_8TH40 U627 ( .A1(n143), .A2(n493), .ZN(n463) );
  AND2V0_8TH40 U628 ( .A1(n494), .A2(n502), .Z(n493) );
  NOR2V0P5_8TH40 U629 ( .A1(inst_i[29]), .A2(inst_i[28]), .ZN(n502) );
  CLKNV1_8TH40 U630 ( .I(n216), .ZN(n195) );
  NOR2V0P5_8TH40 U631 ( .A1(n186), .A2(n193), .ZN(n216) );
  CLKNAND2V1_8TH40 U632 ( .A1(inst_i[27]), .A2(inst_i[26]), .ZN(n193) );
  CLKNV1_8TH40 U633 ( .I(n217), .ZN(n119) );
  AOI21V0_8TH40 U634 ( .A1(n147), .A2(n391), .B(n186), .ZN(n217) );
  NAND3V0P5_8TH40 U635 ( .A1(inst_i[29]), .A2(n494), .A3(inst_i[28]), .ZN(n186) );
  NOR2V0P5_8TH40 U636 ( .A1(inst_i[31]), .A2(inst_i[30]), .ZN(n494) );
  NOR2V0P5_8TH40 U637 ( .A1(n122), .A2(n143), .ZN(n391) );
  NOR2V0P5_8TH40 U638 ( .A1(n497), .A2(inst_i[27]), .ZN(n143) );
  NOR2V0P5_8TH40 U639 ( .A1(inst_i[27]), .A2(inst_i[26]), .ZN(n122) );
  CLKNAND2V1_8TH40 U640 ( .A1(inst_i[27]), .A2(n497), .ZN(n147) );
  CLKNV1_8TH40 U641 ( .I(inst_i[26]), .ZN(n497) );
  CLKNV1_8TH40 U642 ( .I(rst), .ZN(n51) );
endmodule


module gpr ( clk, rst, we, waddr, wdata, re1, raddr1, rdata1, re2, raddr2, 
        rdata2 );
  input [4:0] waddr;
  input [31:0] wdata;
  input [4:0] raddr1;
  output [31:0] rdata1;
  input [4:0] raddr2;
  output [31:0] rdata2;
  input clk, rst, we, re1, re2;
  wire   N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N140, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250;
  wire   [1023:0] regs;

  DQV4_8TH40 regs_reg_3__31_ ( .D(n528), .CK(clk), .Q(regs[927]) );
  DQV4_8TH40 regs_reg_3__30_ ( .D(n527), .CK(clk), .Q(regs[926]) );
  DQV4_8TH40 regs_reg_3__29_ ( .D(n526), .CK(clk), .Q(regs[925]) );
  DQV4_8TH40 regs_reg_3__28_ ( .D(n525), .CK(clk), .Q(regs[924]) );
  DQV4_8TH40 regs_reg_3__27_ ( .D(n524), .CK(clk), .Q(regs[923]) );
  DQV4_8TH40 regs_reg_3__26_ ( .D(n523), .CK(clk), .Q(regs[922]) );
  DQV4_8TH40 regs_reg_3__25_ ( .D(n522), .CK(clk), .Q(regs[921]) );
  DQV4_8TH40 regs_reg_3__24_ ( .D(n521), .CK(clk), .Q(regs[920]) );
  DQV4_8TH40 regs_reg_3__23_ ( .D(n520), .CK(clk), .Q(regs[919]) );
  DQV4_8TH40 regs_reg_3__22_ ( .D(n519), .CK(clk), .Q(regs[918]) );
  DQV4_8TH40 regs_reg_3__21_ ( .D(n518), .CK(clk), .Q(regs[917]) );
  DQV4_8TH40 regs_reg_3__20_ ( .D(n517), .CK(clk), .Q(regs[916]) );
  DQV4_8TH40 regs_reg_3__19_ ( .D(n516), .CK(clk), .Q(regs[915]) );
  DQV4_8TH40 regs_reg_3__18_ ( .D(n515), .CK(clk), .Q(regs[914]) );
  DQV4_8TH40 regs_reg_3__17_ ( .D(n514), .CK(clk), .Q(regs[913]) );
  DQV4_8TH40 regs_reg_3__16_ ( .D(n513), .CK(clk), .Q(regs[912]) );
  DQV4_8TH40 regs_reg_3__15_ ( .D(n512), .CK(clk), .Q(regs[911]) );
  DQV4_8TH40 regs_reg_3__14_ ( .D(n511), .CK(clk), .Q(regs[910]) );
  DQV4_8TH40 regs_reg_3__13_ ( .D(n510), .CK(clk), .Q(regs[909]) );
  DQV4_8TH40 regs_reg_3__12_ ( .D(n509), .CK(clk), .Q(regs[908]) );
  DQV4_8TH40 regs_reg_3__11_ ( .D(n508), .CK(clk), .Q(regs[907]) );
  DQV4_8TH40 regs_reg_3__10_ ( .D(n507), .CK(clk), .Q(regs[906]) );
  DQV4_8TH40 regs_reg_3__9_ ( .D(n506), .CK(clk), .Q(regs[905]) );
  DQV4_8TH40 regs_reg_3__8_ ( .D(n505), .CK(clk), .Q(regs[904]) );
  DQV4_8TH40 regs_reg_3__7_ ( .D(n504), .CK(clk), .Q(regs[903]) );
  DQV4_8TH40 regs_reg_3__6_ ( .D(n503), .CK(clk), .Q(regs[902]) );
  DQV4_8TH40 regs_reg_3__5_ ( .D(n502), .CK(clk), .Q(regs[901]) );
  DQV4_8TH40 regs_reg_3__4_ ( .D(n501), .CK(clk), .Q(regs[900]) );
  DQV4_8TH40 regs_reg_3__3_ ( .D(n500), .CK(clk), .Q(regs[899]) );
  DQV4_8TH40 regs_reg_3__2_ ( .D(n499), .CK(clk), .Q(regs[898]) );
  DQV4_8TH40 regs_reg_3__1_ ( .D(n498), .CK(clk), .Q(regs[897]) );
  DQV4_8TH40 regs_reg_3__0_ ( .D(n497), .CK(clk), .Q(regs[896]) );
  DQV4_8TH40 regs_reg_5__31_ ( .D(n496), .CK(clk), .Q(regs[863]) );
  DQV4_8TH40 regs_reg_5__30_ ( .D(n495), .CK(clk), .Q(regs[862]) );
  DQV4_8TH40 regs_reg_5__29_ ( .D(n494), .CK(clk), .Q(regs[861]) );
  DQV4_8TH40 regs_reg_5__28_ ( .D(n493), .CK(clk), .Q(regs[860]) );
  DQV4_8TH40 regs_reg_5__27_ ( .D(n492), .CK(clk), .Q(regs[859]) );
  DQV4_8TH40 regs_reg_5__26_ ( .D(n491), .CK(clk), .Q(regs[858]) );
  DQV4_8TH40 regs_reg_5__25_ ( .D(n490), .CK(clk), .Q(regs[857]) );
  DQV4_8TH40 regs_reg_5__24_ ( .D(n489), .CK(clk), .Q(regs[856]) );
  DQV4_8TH40 regs_reg_5__23_ ( .D(n488), .CK(clk), .Q(regs[855]) );
  DQV4_8TH40 regs_reg_5__22_ ( .D(n487), .CK(clk), .Q(regs[854]) );
  DQV4_8TH40 regs_reg_5__21_ ( .D(n486), .CK(clk), .Q(regs[853]) );
  DQV4_8TH40 regs_reg_5__20_ ( .D(n485), .CK(clk), .Q(regs[852]) );
  DQV4_8TH40 regs_reg_5__19_ ( .D(n484), .CK(clk), .Q(regs[851]) );
  DQV4_8TH40 regs_reg_5__18_ ( .D(n483), .CK(clk), .Q(regs[850]) );
  DQV4_8TH40 regs_reg_5__17_ ( .D(n482), .CK(clk), .Q(regs[849]) );
  DQV4_8TH40 regs_reg_5__16_ ( .D(n481), .CK(clk), .Q(regs[848]) );
  DQV4_8TH40 regs_reg_5__15_ ( .D(n480), .CK(clk), .Q(regs[847]) );
  DQV4_8TH40 regs_reg_5__14_ ( .D(n479), .CK(clk), .Q(regs[846]) );
  DQV4_8TH40 regs_reg_5__13_ ( .D(n478), .CK(clk), .Q(regs[845]) );
  DQV4_8TH40 regs_reg_5__12_ ( .D(n477), .CK(clk), .Q(regs[844]) );
  DQV4_8TH40 regs_reg_5__11_ ( .D(n476), .CK(clk), .Q(regs[843]) );
  DQV4_8TH40 regs_reg_5__10_ ( .D(n475), .CK(clk), .Q(regs[842]) );
  DQV4_8TH40 regs_reg_5__9_ ( .D(n474), .CK(clk), .Q(regs[841]) );
  DQV4_8TH40 regs_reg_5__8_ ( .D(n473), .CK(clk), .Q(regs[840]) );
  DQV4_8TH40 regs_reg_5__7_ ( .D(n472), .CK(clk), .Q(regs[839]) );
  DQV4_8TH40 regs_reg_5__6_ ( .D(n471), .CK(clk), .Q(regs[838]) );
  DQV4_8TH40 regs_reg_5__5_ ( .D(n470), .CK(clk), .Q(regs[837]) );
  DQV4_8TH40 regs_reg_5__4_ ( .D(n469), .CK(clk), .Q(regs[836]) );
  DQV4_8TH40 regs_reg_5__3_ ( .D(n468), .CK(clk), .Q(regs[835]) );
  DQV4_8TH40 regs_reg_5__2_ ( .D(n467), .CK(clk), .Q(regs[834]) );
  DQV4_8TH40 regs_reg_5__1_ ( .D(n466), .CK(clk), .Q(regs[833]) );
  DQV4_8TH40 regs_reg_5__0_ ( .D(n465), .CK(clk), .Q(regs[832]) );
  DQV4_8TH40 regs_reg_6__31_ ( .D(n464), .CK(clk), .Q(regs[831]) );
  DQV4_8TH40 regs_reg_6__30_ ( .D(n463), .CK(clk), .Q(regs[830]) );
  DQV4_8TH40 regs_reg_6__29_ ( .D(n462), .CK(clk), .Q(regs[829]) );
  DQV4_8TH40 regs_reg_6__28_ ( .D(n461), .CK(clk), .Q(regs[828]) );
  DQV4_8TH40 regs_reg_6__27_ ( .D(n460), .CK(clk), .Q(regs[827]) );
  DQV4_8TH40 regs_reg_6__26_ ( .D(n459), .CK(clk), .Q(regs[826]) );
  DQV4_8TH40 regs_reg_6__25_ ( .D(n458), .CK(clk), .Q(regs[825]) );
  DQV4_8TH40 regs_reg_6__24_ ( .D(n457), .CK(clk), .Q(regs[824]) );
  DQV4_8TH40 regs_reg_6__23_ ( .D(n456), .CK(clk), .Q(regs[823]) );
  DQV4_8TH40 regs_reg_6__22_ ( .D(n455), .CK(clk), .Q(regs[822]) );
  DQV4_8TH40 regs_reg_6__21_ ( .D(n454), .CK(clk), .Q(regs[821]) );
  DQV4_8TH40 regs_reg_6__20_ ( .D(n453), .CK(clk), .Q(regs[820]) );
  DQV4_8TH40 regs_reg_6__19_ ( .D(n452), .CK(clk), .Q(regs[819]) );
  DQV4_8TH40 regs_reg_6__18_ ( .D(n451), .CK(clk), .Q(regs[818]) );
  DQV4_8TH40 regs_reg_6__17_ ( .D(n450), .CK(clk), .Q(regs[817]) );
  DQV4_8TH40 regs_reg_6__16_ ( .D(n449), .CK(clk), .Q(regs[816]) );
  DQV4_8TH40 regs_reg_6__15_ ( .D(n448), .CK(clk), .Q(regs[815]) );
  DQV4_8TH40 regs_reg_6__14_ ( .D(n447), .CK(clk), .Q(regs[814]) );
  DQV4_8TH40 regs_reg_6__13_ ( .D(n446), .CK(clk), .Q(regs[813]) );
  DQV4_8TH40 regs_reg_6__12_ ( .D(n445), .CK(clk), .Q(regs[812]) );
  DQV4_8TH40 regs_reg_6__11_ ( .D(n444), .CK(clk), .Q(regs[811]) );
  DQV4_8TH40 regs_reg_6__10_ ( .D(n443), .CK(clk), .Q(regs[810]) );
  DQV4_8TH40 regs_reg_6__9_ ( .D(n442), .CK(clk), .Q(regs[809]) );
  DQV4_8TH40 regs_reg_6__8_ ( .D(n441), .CK(clk), .Q(regs[808]) );
  DQV4_8TH40 regs_reg_6__7_ ( .D(n440), .CK(clk), .Q(regs[807]) );
  DQV4_8TH40 regs_reg_6__6_ ( .D(n439), .CK(clk), .Q(regs[806]) );
  DQV4_8TH40 regs_reg_6__5_ ( .D(n438), .CK(clk), .Q(regs[805]) );
  DQV4_8TH40 regs_reg_6__4_ ( .D(n437), .CK(clk), .Q(regs[804]) );
  DQV4_8TH40 regs_reg_6__3_ ( .D(n436), .CK(clk), .Q(regs[803]) );
  DQV4_8TH40 regs_reg_6__2_ ( .D(n435), .CK(clk), .Q(regs[802]) );
  DQV4_8TH40 regs_reg_6__1_ ( .D(n434), .CK(clk), .Q(regs[801]) );
  DQV4_8TH40 regs_reg_6__0_ ( .D(n433), .CK(clk), .Q(regs[800]) );
  DQV4_8TH40 regs_reg_7__31_ ( .D(n432), .CK(clk), .Q(regs[799]) );
  DQV4_8TH40 regs_reg_7__30_ ( .D(n431), .CK(clk), .Q(regs[798]) );
  DQV4_8TH40 regs_reg_7__29_ ( .D(n430), .CK(clk), .Q(regs[797]) );
  DQV4_8TH40 regs_reg_7__28_ ( .D(n429), .CK(clk), .Q(regs[796]) );
  DQV4_8TH40 regs_reg_7__27_ ( .D(n428), .CK(clk), .Q(regs[795]) );
  DQV4_8TH40 regs_reg_7__26_ ( .D(n427), .CK(clk), .Q(regs[794]) );
  DQV4_8TH40 regs_reg_7__25_ ( .D(n426), .CK(clk), .Q(regs[793]) );
  DQV4_8TH40 regs_reg_7__24_ ( .D(n425), .CK(clk), .Q(regs[792]) );
  DQV4_8TH40 regs_reg_7__23_ ( .D(n424), .CK(clk), .Q(regs[791]) );
  DQV4_8TH40 regs_reg_7__22_ ( .D(n423), .CK(clk), .Q(regs[790]) );
  DQV4_8TH40 regs_reg_7__21_ ( .D(n422), .CK(clk), .Q(regs[789]) );
  DQV4_8TH40 regs_reg_7__20_ ( .D(n421), .CK(clk), .Q(regs[788]) );
  DQV4_8TH40 regs_reg_7__19_ ( .D(n420), .CK(clk), .Q(regs[787]) );
  DQV4_8TH40 regs_reg_7__18_ ( .D(n419), .CK(clk), .Q(regs[786]) );
  DQV4_8TH40 regs_reg_7__17_ ( .D(n418), .CK(clk), .Q(regs[785]) );
  DQV4_8TH40 regs_reg_7__16_ ( .D(n417), .CK(clk), .Q(regs[784]) );
  DQV4_8TH40 regs_reg_7__15_ ( .D(n416), .CK(clk), .Q(regs[783]) );
  DQV4_8TH40 regs_reg_7__14_ ( .D(n415), .CK(clk), .Q(regs[782]) );
  DQV4_8TH40 regs_reg_7__13_ ( .D(n414), .CK(clk), .Q(regs[781]) );
  DQV4_8TH40 regs_reg_7__12_ ( .D(n413), .CK(clk), .Q(regs[780]) );
  DQV4_8TH40 regs_reg_7__11_ ( .D(n412), .CK(clk), .Q(regs[779]) );
  DQV4_8TH40 regs_reg_7__10_ ( .D(n411), .CK(clk), .Q(regs[778]) );
  DQV4_8TH40 regs_reg_7__9_ ( .D(n410), .CK(clk), .Q(regs[777]) );
  DQV4_8TH40 regs_reg_7__8_ ( .D(n409), .CK(clk), .Q(regs[776]) );
  DQV4_8TH40 regs_reg_7__7_ ( .D(n408), .CK(clk), .Q(regs[775]) );
  DQV4_8TH40 regs_reg_7__6_ ( .D(n407), .CK(clk), .Q(regs[774]) );
  DQV4_8TH40 regs_reg_7__5_ ( .D(n406), .CK(clk), .Q(regs[773]) );
  DQV4_8TH40 regs_reg_7__4_ ( .D(n405), .CK(clk), .Q(regs[772]) );
  DQV4_8TH40 regs_reg_7__3_ ( .D(n404), .CK(clk), .Q(regs[771]) );
  DQV4_8TH40 regs_reg_7__2_ ( .D(n403), .CK(clk), .Q(regs[770]) );
  DQV4_8TH40 regs_reg_7__1_ ( .D(n402), .CK(clk), .Q(regs[769]) );
  DQV4_8TH40 regs_reg_7__0_ ( .D(n401), .CK(clk), .Q(regs[768]) );
  DQV4_8TH40 regs_reg_11__31_ ( .D(n400), .CK(clk), .Q(regs[671]) );
  DQV4_8TH40 regs_reg_11__30_ ( .D(n399), .CK(clk), .Q(regs[670]) );
  DQV4_8TH40 regs_reg_11__29_ ( .D(n398), .CK(clk), .Q(regs[669]) );
  DQV4_8TH40 regs_reg_11__28_ ( .D(n397), .CK(clk), .Q(regs[668]) );
  DQV4_8TH40 regs_reg_11__27_ ( .D(n396), .CK(clk), .Q(regs[667]) );
  DQV4_8TH40 regs_reg_11__26_ ( .D(n395), .CK(clk), .Q(regs[666]) );
  DQV4_8TH40 regs_reg_11__25_ ( .D(n394), .CK(clk), .Q(regs[665]) );
  DQV4_8TH40 regs_reg_11__24_ ( .D(n393), .CK(clk), .Q(regs[664]) );
  DQV4_8TH40 regs_reg_11__23_ ( .D(n392), .CK(clk), .Q(regs[663]) );
  DQV4_8TH40 regs_reg_11__22_ ( .D(n391), .CK(clk), .Q(regs[662]) );
  DQV4_8TH40 regs_reg_11__21_ ( .D(n390), .CK(clk), .Q(regs[661]) );
  DQV4_8TH40 regs_reg_11__20_ ( .D(n389), .CK(clk), .Q(regs[660]) );
  DQV4_8TH40 regs_reg_11__19_ ( .D(n388), .CK(clk), .Q(regs[659]) );
  DQV4_8TH40 regs_reg_11__18_ ( .D(n387), .CK(clk), .Q(regs[658]) );
  DQV4_8TH40 regs_reg_11__17_ ( .D(n386), .CK(clk), .Q(regs[657]) );
  DQV4_8TH40 regs_reg_11__16_ ( .D(n385), .CK(clk), .Q(regs[656]) );
  DQV4_8TH40 regs_reg_11__15_ ( .D(n384), .CK(clk), .Q(regs[655]) );
  DQV4_8TH40 regs_reg_11__14_ ( .D(n383), .CK(clk), .Q(regs[654]) );
  DQV4_8TH40 regs_reg_11__13_ ( .D(n382), .CK(clk), .Q(regs[653]) );
  DQV4_8TH40 regs_reg_11__12_ ( .D(n381), .CK(clk), .Q(regs[652]) );
  DQV4_8TH40 regs_reg_11__11_ ( .D(n380), .CK(clk), .Q(regs[651]) );
  DQV4_8TH40 regs_reg_11__10_ ( .D(n379), .CK(clk), .Q(regs[650]) );
  DQV4_8TH40 regs_reg_11__9_ ( .D(n378), .CK(clk), .Q(regs[649]) );
  DQV4_8TH40 regs_reg_11__8_ ( .D(n377), .CK(clk), .Q(regs[648]) );
  DQV4_8TH40 regs_reg_11__7_ ( .D(n376), .CK(clk), .Q(regs[647]) );
  DQV4_8TH40 regs_reg_11__6_ ( .D(n375), .CK(clk), .Q(regs[646]) );
  DQV4_8TH40 regs_reg_11__5_ ( .D(n374), .CK(clk), .Q(regs[645]) );
  DQV4_8TH40 regs_reg_11__4_ ( .D(n373), .CK(clk), .Q(regs[644]) );
  DQV4_8TH40 regs_reg_11__3_ ( .D(n372), .CK(clk), .Q(regs[643]) );
  DQV4_8TH40 regs_reg_11__2_ ( .D(n371), .CK(clk), .Q(regs[642]) );
  DQV4_8TH40 regs_reg_11__1_ ( .D(n370), .CK(clk), .Q(regs[641]) );
  DQV4_8TH40 regs_reg_11__0_ ( .D(n369), .CK(clk), .Q(regs[640]) );
  DQV4_8TH40 regs_reg_13__31_ ( .D(n368), .CK(clk), .Q(regs[607]) );
  DQV4_8TH40 regs_reg_13__30_ ( .D(n367), .CK(clk), .Q(regs[606]) );
  DQV4_8TH40 regs_reg_13__29_ ( .D(n366), .CK(clk), .Q(regs[605]) );
  DQV4_8TH40 regs_reg_13__28_ ( .D(n365), .CK(clk), .Q(regs[604]) );
  DQV4_8TH40 regs_reg_13__27_ ( .D(n364), .CK(clk), .Q(regs[603]) );
  DQV4_8TH40 regs_reg_13__26_ ( .D(n363), .CK(clk), .Q(regs[602]) );
  DQV4_8TH40 regs_reg_13__25_ ( .D(n362), .CK(clk), .Q(regs[601]) );
  DQV4_8TH40 regs_reg_13__24_ ( .D(n361), .CK(clk), .Q(regs[600]) );
  DQV4_8TH40 regs_reg_13__23_ ( .D(n360), .CK(clk), .Q(regs[599]) );
  DQV4_8TH40 regs_reg_13__22_ ( .D(n359), .CK(clk), .Q(regs[598]) );
  DQV4_8TH40 regs_reg_13__21_ ( .D(n358), .CK(clk), .Q(regs[597]) );
  DQV4_8TH40 regs_reg_13__20_ ( .D(n357), .CK(clk), .Q(regs[596]) );
  DQV4_8TH40 regs_reg_13__19_ ( .D(n356), .CK(clk), .Q(regs[595]) );
  DQV4_8TH40 regs_reg_13__18_ ( .D(n355), .CK(clk), .Q(regs[594]) );
  DQV4_8TH40 regs_reg_13__17_ ( .D(n354), .CK(clk), .Q(regs[593]) );
  DQV4_8TH40 regs_reg_13__16_ ( .D(n353), .CK(clk), .Q(regs[592]) );
  DQV4_8TH40 regs_reg_13__15_ ( .D(n352), .CK(clk), .Q(regs[591]) );
  DQV4_8TH40 regs_reg_13__14_ ( .D(n351), .CK(clk), .Q(regs[590]) );
  DQV4_8TH40 regs_reg_13__13_ ( .D(n350), .CK(clk), .Q(regs[589]) );
  DQV4_8TH40 regs_reg_13__12_ ( .D(n349), .CK(clk), .Q(regs[588]) );
  DQV4_8TH40 regs_reg_13__11_ ( .D(n348), .CK(clk), .Q(regs[587]) );
  DQV4_8TH40 regs_reg_13__10_ ( .D(n347), .CK(clk), .Q(regs[586]) );
  DQV4_8TH40 regs_reg_13__9_ ( .D(n346), .CK(clk), .Q(regs[585]) );
  DQV4_8TH40 regs_reg_13__8_ ( .D(n345), .CK(clk), .Q(regs[584]) );
  DQV4_8TH40 regs_reg_13__7_ ( .D(n344), .CK(clk), .Q(regs[583]) );
  DQV4_8TH40 regs_reg_13__6_ ( .D(n343), .CK(clk), .Q(regs[582]) );
  DQV4_8TH40 regs_reg_13__5_ ( .D(n342), .CK(clk), .Q(regs[581]) );
  DQV4_8TH40 regs_reg_13__4_ ( .D(n341), .CK(clk), .Q(regs[580]) );
  DQV4_8TH40 regs_reg_13__3_ ( .D(n340), .CK(clk), .Q(regs[579]) );
  DQV4_8TH40 regs_reg_13__2_ ( .D(n339), .CK(clk), .Q(regs[578]) );
  DQV4_8TH40 regs_reg_13__1_ ( .D(n338), .CK(clk), .Q(regs[577]) );
  DQV4_8TH40 regs_reg_13__0_ ( .D(n337), .CK(clk), .Q(regs[576]) );
  DQV4_8TH40 regs_reg_14__31_ ( .D(n336), .CK(clk), .Q(regs[575]) );
  DQV4_8TH40 regs_reg_14__30_ ( .D(n335), .CK(clk), .Q(regs[574]) );
  DQV4_8TH40 regs_reg_14__29_ ( .D(n334), .CK(clk), .Q(regs[573]) );
  DQV4_8TH40 regs_reg_14__28_ ( .D(n333), .CK(clk), .Q(regs[572]) );
  DQV4_8TH40 regs_reg_14__27_ ( .D(n332), .CK(clk), .Q(regs[571]) );
  DQV4_8TH40 regs_reg_14__26_ ( .D(n331), .CK(clk), .Q(regs[570]) );
  DQV4_8TH40 regs_reg_14__25_ ( .D(n330), .CK(clk), .Q(regs[569]) );
  DQV4_8TH40 regs_reg_14__24_ ( .D(n329), .CK(clk), .Q(regs[568]) );
  DQV4_8TH40 regs_reg_14__23_ ( .D(n328), .CK(clk), .Q(regs[567]) );
  DQV4_8TH40 regs_reg_14__22_ ( .D(n327), .CK(clk), .Q(regs[566]) );
  DQV4_8TH40 regs_reg_14__21_ ( .D(n326), .CK(clk), .Q(regs[565]) );
  DQV4_8TH40 regs_reg_14__20_ ( .D(n325), .CK(clk), .Q(regs[564]) );
  DQV4_8TH40 regs_reg_14__19_ ( .D(n324), .CK(clk), .Q(regs[563]) );
  DQV4_8TH40 regs_reg_14__18_ ( .D(n323), .CK(clk), .Q(regs[562]) );
  DQV4_8TH40 regs_reg_14__17_ ( .D(n322), .CK(clk), .Q(regs[561]) );
  DQV4_8TH40 regs_reg_14__16_ ( .D(n321), .CK(clk), .Q(regs[560]) );
  DQV4_8TH40 regs_reg_14__15_ ( .D(n320), .CK(clk), .Q(regs[559]) );
  DQV4_8TH40 regs_reg_14__14_ ( .D(n319), .CK(clk), .Q(regs[558]) );
  DQV4_8TH40 regs_reg_14__13_ ( .D(n318), .CK(clk), .Q(regs[557]) );
  DQV4_8TH40 regs_reg_14__12_ ( .D(n317), .CK(clk), .Q(regs[556]) );
  DQV4_8TH40 regs_reg_14__11_ ( .D(n316), .CK(clk), .Q(regs[555]) );
  DQV4_8TH40 regs_reg_14__10_ ( .D(n315), .CK(clk), .Q(regs[554]) );
  DQV4_8TH40 regs_reg_14__9_ ( .D(n314), .CK(clk), .Q(regs[553]) );
  DQV4_8TH40 regs_reg_14__8_ ( .D(n313), .CK(clk), .Q(regs[552]) );
  DQV4_8TH40 regs_reg_14__7_ ( .D(n312), .CK(clk), .Q(regs[551]) );
  DQV4_8TH40 regs_reg_14__6_ ( .D(n311), .CK(clk), .Q(regs[550]) );
  DQV4_8TH40 regs_reg_14__5_ ( .D(n310), .CK(clk), .Q(regs[549]) );
  DQV4_8TH40 regs_reg_14__4_ ( .D(n309), .CK(clk), .Q(regs[548]) );
  DQV4_8TH40 regs_reg_14__3_ ( .D(n308), .CK(clk), .Q(regs[547]) );
  DQV4_8TH40 regs_reg_14__2_ ( .D(n307), .CK(clk), .Q(regs[546]) );
  DQV4_8TH40 regs_reg_14__1_ ( .D(n306), .CK(clk), .Q(regs[545]) );
  DQV4_8TH40 regs_reg_14__0_ ( .D(n305), .CK(clk), .Q(regs[544]) );
  DQV4_8TH40 regs_reg_15__31_ ( .D(n304), .CK(clk), .Q(regs[543]) );
  DQV4_8TH40 regs_reg_15__30_ ( .D(n303), .CK(clk), .Q(regs[542]) );
  DQV4_8TH40 regs_reg_15__29_ ( .D(n302), .CK(clk), .Q(regs[541]) );
  DQV4_8TH40 regs_reg_15__28_ ( .D(n301), .CK(clk), .Q(regs[540]) );
  DQV4_8TH40 regs_reg_15__27_ ( .D(n300), .CK(clk), .Q(regs[539]) );
  DQV4_8TH40 regs_reg_15__26_ ( .D(n299), .CK(clk), .Q(regs[538]) );
  DQV4_8TH40 regs_reg_15__25_ ( .D(n298), .CK(clk), .Q(regs[537]) );
  DQV4_8TH40 regs_reg_15__24_ ( .D(n297), .CK(clk), .Q(regs[536]) );
  DQV4_8TH40 regs_reg_15__23_ ( .D(n296), .CK(clk), .Q(regs[535]) );
  DQV4_8TH40 regs_reg_15__22_ ( .D(n295), .CK(clk), .Q(regs[534]) );
  DQV4_8TH40 regs_reg_15__21_ ( .D(n294), .CK(clk), .Q(regs[533]) );
  DQV4_8TH40 regs_reg_15__20_ ( .D(n293), .CK(clk), .Q(regs[532]) );
  DQV4_8TH40 regs_reg_15__19_ ( .D(n292), .CK(clk), .Q(regs[531]) );
  DQV4_8TH40 regs_reg_15__18_ ( .D(n291), .CK(clk), .Q(regs[530]) );
  DQV4_8TH40 regs_reg_15__17_ ( .D(n290), .CK(clk), .Q(regs[529]) );
  DQV4_8TH40 regs_reg_15__16_ ( .D(n289), .CK(clk), .Q(regs[528]) );
  DQV4_8TH40 regs_reg_15__15_ ( .D(n288), .CK(clk), .Q(regs[527]) );
  DQV4_8TH40 regs_reg_15__14_ ( .D(n287), .CK(clk), .Q(regs[526]) );
  DQV4_8TH40 regs_reg_15__13_ ( .D(n286), .CK(clk), .Q(regs[525]) );
  DQV4_8TH40 regs_reg_15__12_ ( .D(n285), .CK(clk), .Q(regs[524]) );
  DQV4_8TH40 regs_reg_15__11_ ( .D(n284), .CK(clk), .Q(regs[523]) );
  DQV4_8TH40 regs_reg_15__10_ ( .D(n283), .CK(clk), .Q(regs[522]) );
  DQV4_8TH40 regs_reg_15__9_ ( .D(n282), .CK(clk), .Q(regs[521]) );
  DQV4_8TH40 regs_reg_15__8_ ( .D(n281), .CK(clk), .Q(regs[520]) );
  DQV4_8TH40 regs_reg_15__7_ ( .D(n280), .CK(clk), .Q(regs[519]) );
  DQV4_8TH40 regs_reg_15__6_ ( .D(n279), .CK(clk), .Q(regs[518]) );
  DQV4_8TH40 regs_reg_15__5_ ( .D(n278), .CK(clk), .Q(regs[517]) );
  DQV4_8TH40 regs_reg_15__4_ ( .D(n277), .CK(clk), .Q(regs[516]) );
  DQV4_8TH40 regs_reg_15__3_ ( .D(n276), .CK(clk), .Q(regs[515]) );
  DQV4_8TH40 regs_reg_15__2_ ( .D(n275), .CK(clk), .Q(regs[514]) );
  DQV4_8TH40 regs_reg_15__1_ ( .D(n274), .CK(clk), .Q(regs[513]) );
  DQV4_8TH40 regs_reg_15__0_ ( .D(n273), .CK(clk), .Q(regs[512]) );
  DQV4_8TH40 regs_reg_23__31_ ( .D(n272), .CK(clk), .Q(regs[287]) );
  DQV4_8TH40 regs_reg_23__30_ ( .D(n271), .CK(clk), .Q(regs[286]) );
  DQV4_8TH40 regs_reg_23__29_ ( .D(n270), .CK(clk), .Q(regs[285]) );
  DQV4_8TH40 regs_reg_23__28_ ( .D(n269), .CK(clk), .Q(regs[284]) );
  DQV4_8TH40 regs_reg_23__27_ ( .D(n268), .CK(clk), .Q(regs[283]) );
  DQV4_8TH40 regs_reg_23__26_ ( .D(n267), .CK(clk), .Q(regs[282]) );
  DQV4_8TH40 regs_reg_23__25_ ( .D(n266), .CK(clk), .Q(regs[281]) );
  DQV4_8TH40 regs_reg_23__24_ ( .D(n265), .CK(clk), .Q(regs[280]) );
  DQV4_8TH40 regs_reg_23__23_ ( .D(n264), .CK(clk), .Q(regs[279]) );
  DQV4_8TH40 regs_reg_23__22_ ( .D(n263), .CK(clk), .Q(regs[278]) );
  DQV4_8TH40 regs_reg_23__21_ ( .D(n262), .CK(clk), .Q(regs[277]) );
  DQV4_8TH40 regs_reg_23__20_ ( .D(n261), .CK(clk), .Q(regs[276]) );
  DQV4_8TH40 regs_reg_23__19_ ( .D(n260), .CK(clk), .Q(regs[275]) );
  DQV4_8TH40 regs_reg_23__18_ ( .D(n259), .CK(clk), .Q(regs[274]) );
  DQV4_8TH40 regs_reg_23__17_ ( .D(n258), .CK(clk), .Q(regs[273]) );
  DQV4_8TH40 regs_reg_23__16_ ( .D(n257), .CK(clk), .Q(regs[272]) );
  DQV4_8TH40 regs_reg_23__15_ ( .D(n256), .CK(clk), .Q(regs[271]) );
  DQV4_8TH40 regs_reg_23__14_ ( .D(n255), .CK(clk), .Q(regs[270]) );
  DQV4_8TH40 regs_reg_23__13_ ( .D(n254), .CK(clk), .Q(regs[269]) );
  DQV4_8TH40 regs_reg_23__12_ ( .D(n253), .CK(clk), .Q(regs[268]) );
  DQV4_8TH40 regs_reg_23__11_ ( .D(n252), .CK(clk), .Q(regs[267]) );
  DQV4_8TH40 regs_reg_23__10_ ( .D(n251), .CK(clk), .Q(regs[266]) );
  DQV4_8TH40 regs_reg_23__9_ ( .D(n250), .CK(clk), .Q(regs[265]) );
  DQV4_8TH40 regs_reg_23__8_ ( .D(n249), .CK(clk), .Q(regs[264]) );
  DQV4_8TH40 regs_reg_23__7_ ( .D(n248), .CK(clk), .Q(regs[263]) );
  DQV4_8TH40 regs_reg_23__6_ ( .D(n247), .CK(clk), .Q(regs[262]) );
  DQV4_8TH40 regs_reg_23__5_ ( .D(n246), .CK(clk), .Q(regs[261]) );
  DQV4_8TH40 regs_reg_23__4_ ( .D(n245), .CK(clk), .Q(regs[260]) );
  DQV4_8TH40 regs_reg_23__3_ ( .D(n244), .CK(clk), .Q(regs[259]) );
  DQV4_8TH40 regs_reg_23__2_ ( .D(n243), .CK(clk), .Q(regs[258]) );
  DQV4_8TH40 regs_reg_23__1_ ( .D(n242), .CK(clk), .Q(regs[257]) );
  DQV4_8TH40 regs_reg_23__0_ ( .D(n241), .CK(clk), .Q(regs[256]) );
  DQV4_8TH40 regs_reg_27__31_ ( .D(n240), .CK(clk), .Q(regs[159]) );
  DQV4_8TH40 regs_reg_27__30_ ( .D(n239), .CK(clk), .Q(regs[158]) );
  DQV4_8TH40 regs_reg_27__29_ ( .D(n238), .CK(clk), .Q(regs[157]) );
  DQV4_8TH40 regs_reg_27__28_ ( .D(n237), .CK(clk), .Q(regs[156]) );
  DQV4_8TH40 regs_reg_27__27_ ( .D(n236), .CK(clk), .Q(regs[155]) );
  DQV4_8TH40 regs_reg_27__26_ ( .D(n235), .CK(clk), .Q(regs[154]) );
  DQV4_8TH40 regs_reg_27__25_ ( .D(n234), .CK(clk), .Q(regs[153]) );
  DQV4_8TH40 regs_reg_27__24_ ( .D(n233), .CK(clk), .Q(regs[152]) );
  DQV4_8TH40 regs_reg_27__23_ ( .D(n232), .CK(clk), .Q(regs[151]) );
  DQV4_8TH40 regs_reg_27__22_ ( .D(n231), .CK(clk), .Q(regs[150]) );
  DQV4_8TH40 regs_reg_27__21_ ( .D(n230), .CK(clk), .Q(regs[149]) );
  DQV4_8TH40 regs_reg_27__20_ ( .D(n229), .CK(clk), .Q(regs[148]) );
  DQV4_8TH40 regs_reg_27__19_ ( .D(n228), .CK(clk), .Q(regs[147]) );
  DQV4_8TH40 regs_reg_27__18_ ( .D(n227), .CK(clk), .Q(regs[146]) );
  DQV4_8TH40 regs_reg_27__17_ ( .D(n226), .CK(clk), .Q(regs[145]) );
  DQV4_8TH40 regs_reg_27__16_ ( .D(n225), .CK(clk), .Q(regs[144]) );
  DQV4_8TH40 regs_reg_27__15_ ( .D(n224), .CK(clk), .Q(regs[143]) );
  DQV4_8TH40 regs_reg_27__14_ ( .D(n223), .CK(clk), .Q(regs[142]) );
  DQV4_8TH40 regs_reg_27__13_ ( .D(n222), .CK(clk), .Q(regs[141]) );
  DQV4_8TH40 regs_reg_27__12_ ( .D(n221), .CK(clk), .Q(regs[140]) );
  DQV4_8TH40 regs_reg_27__11_ ( .D(n220), .CK(clk), .Q(regs[139]) );
  DQV4_8TH40 regs_reg_27__10_ ( .D(n219), .CK(clk), .Q(regs[138]) );
  DQV4_8TH40 regs_reg_27__9_ ( .D(n218), .CK(clk), .Q(regs[137]) );
  DQV4_8TH40 regs_reg_27__8_ ( .D(n217), .CK(clk), .Q(regs[136]) );
  DQV4_8TH40 regs_reg_27__7_ ( .D(n216), .CK(clk), .Q(regs[135]) );
  DQV4_8TH40 regs_reg_27__6_ ( .D(n215), .CK(clk), .Q(regs[134]) );
  DQV4_8TH40 regs_reg_27__5_ ( .D(n214), .CK(clk), .Q(regs[133]) );
  DQV4_8TH40 regs_reg_27__4_ ( .D(n213), .CK(clk), .Q(regs[132]) );
  DQV4_8TH40 regs_reg_27__3_ ( .D(n212), .CK(clk), .Q(regs[131]) );
  DQV4_8TH40 regs_reg_27__2_ ( .D(n211), .CK(clk), .Q(regs[130]) );
  DQV4_8TH40 regs_reg_27__1_ ( .D(n210), .CK(clk), .Q(regs[129]) );
  DQV4_8TH40 regs_reg_27__0_ ( .D(n209), .CK(clk), .Q(regs[128]) );
  DQV4_8TH40 regs_reg_29__31_ ( .D(n208), .CK(clk), .Q(regs[95]) );
  DQV4_8TH40 regs_reg_29__30_ ( .D(n207), .CK(clk), .Q(regs[94]) );
  DQV4_8TH40 regs_reg_29__29_ ( .D(n206), .CK(clk), .Q(regs[93]) );
  DQV4_8TH40 regs_reg_29__28_ ( .D(n205), .CK(clk), .Q(regs[92]) );
  DQV4_8TH40 regs_reg_29__27_ ( .D(n204), .CK(clk), .Q(regs[91]) );
  DQV4_8TH40 regs_reg_29__26_ ( .D(n203), .CK(clk), .Q(regs[90]) );
  DQV4_8TH40 regs_reg_29__25_ ( .D(n202), .CK(clk), .Q(regs[89]) );
  DQV4_8TH40 regs_reg_29__24_ ( .D(n201), .CK(clk), .Q(regs[88]) );
  DQV4_8TH40 regs_reg_29__23_ ( .D(n200), .CK(clk), .Q(regs[87]) );
  DQV4_8TH40 regs_reg_29__22_ ( .D(n199), .CK(clk), .Q(regs[86]) );
  DQV4_8TH40 regs_reg_29__21_ ( .D(n198), .CK(clk), .Q(regs[85]) );
  DQV4_8TH40 regs_reg_29__20_ ( .D(n197), .CK(clk), .Q(regs[84]) );
  DQV4_8TH40 regs_reg_29__19_ ( .D(n196), .CK(clk), .Q(regs[83]) );
  DQV4_8TH40 regs_reg_29__18_ ( .D(n195), .CK(clk), .Q(regs[82]) );
  DQV4_8TH40 regs_reg_29__17_ ( .D(n194), .CK(clk), .Q(regs[81]) );
  DQV4_8TH40 regs_reg_29__16_ ( .D(n193), .CK(clk), .Q(regs[80]) );
  DQV4_8TH40 regs_reg_29__15_ ( .D(n192), .CK(clk), .Q(regs[79]) );
  DQV4_8TH40 regs_reg_29__14_ ( .D(n191), .CK(clk), .Q(regs[78]) );
  DQV4_8TH40 regs_reg_29__13_ ( .D(n190), .CK(clk), .Q(regs[77]) );
  DQV4_8TH40 regs_reg_29__12_ ( .D(n189), .CK(clk), .Q(regs[76]) );
  DQV4_8TH40 regs_reg_29__11_ ( .D(n188), .CK(clk), .Q(regs[75]) );
  DQV4_8TH40 regs_reg_29__10_ ( .D(n187), .CK(clk), .Q(regs[74]) );
  DQV4_8TH40 regs_reg_29__9_ ( .D(n186), .CK(clk), .Q(regs[73]) );
  DQV4_8TH40 regs_reg_29__8_ ( .D(n185), .CK(clk), .Q(regs[72]) );
  DQV4_8TH40 regs_reg_29__7_ ( .D(n184), .CK(clk), .Q(regs[71]) );
  DQV4_8TH40 regs_reg_29__6_ ( .D(n183), .CK(clk), .Q(regs[70]) );
  DQV4_8TH40 regs_reg_29__5_ ( .D(n182), .CK(clk), .Q(regs[69]) );
  DQV4_8TH40 regs_reg_29__4_ ( .D(n181), .CK(clk), .Q(regs[68]) );
  DQV4_8TH40 regs_reg_29__3_ ( .D(n180), .CK(clk), .Q(regs[67]) );
  DQV4_8TH40 regs_reg_29__2_ ( .D(n179), .CK(clk), .Q(regs[66]) );
  DQV4_8TH40 regs_reg_29__1_ ( .D(n178), .CK(clk), .Q(regs[65]) );
  DQV4_8TH40 regs_reg_29__0_ ( .D(n177), .CK(clk), .Q(regs[64]) );
  DQV4_8TH40 regs_reg_30__31_ ( .D(n176), .CK(clk), .Q(regs[63]) );
  DQV4_8TH40 regs_reg_30__30_ ( .D(n175), .CK(clk), .Q(regs[62]) );
  DQV4_8TH40 regs_reg_30__29_ ( .D(n174), .CK(clk), .Q(regs[61]) );
  DQV4_8TH40 regs_reg_30__28_ ( .D(n173), .CK(clk), .Q(regs[60]) );
  DQV4_8TH40 regs_reg_30__27_ ( .D(n172), .CK(clk), .Q(regs[59]) );
  DQV4_8TH40 regs_reg_30__26_ ( .D(n171), .CK(clk), .Q(regs[58]) );
  DQV4_8TH40 regs_reg_30__25_ ( .D(n170), .CK(clk), .Q(regs[57]) );
  DQV4_8TH40 regs_reg_30__24_ ( .D(n169), .CK(clk), .Q(regs[56]) );
  DQV4_8TH40 regs_reg_30__23_ ( .D(n168), .CK(clk), .Q(regs[55]) );
  DQV4_8TH40 regs_reg_30__22_ ( .D(n167), .CK(clk), .Q(regs[54]) );
  DQV4_8TH40 regs_reg_30__21_ ( .D(n166), .CK(clk), .Q(regs[53]) );
  DQV4_8TH40 regs_reg_30__20_ ( .D(n165), .CK(clk), .Q(regs[52]) );
  DQV4_8TH40 regs_reg_30__19_ ( .D(n164), .CK(clk), .Q(regs[51]) );
  DQV4_8TH40 regs_reg_30__18_ ( .D(n163), .CK(clk), .Q(regs[50]) );
  DQV4_8TH40 regs_reg_30__17_ ( .D(n162), .CK(clk), .Q(regs[49]) );
  DQV4_8TH40 regs_reg_30__16_ ( .D(n161), .CK(clk), .Q(regs[48]) );
  DQV4_8TH40 regs_reg_30__15_ ( .D(n160), .CK(clk), .Q(regs[47]) );
  DQV4_8TH40 regs_reg_30__14_ ( .D(n159), .CK(clk), .Q(regs[46]) );
  DQV4_8TH40 regs_reg_30__13_ ( .D(n158), .CK(clk), .Q(regs[45]) );
  DQV4_8TH40 regs_reg_30__12_ ( .D(n157), .CK(clk), .Q(regs[44]) );
  DQV4_8TH40 regs_reg_30__11_ ( .D(n156), .CK(clk), .Q(regs[43]) );
  DQV4_8TH40 regs_reg_30__10_ ( .D(n155), .CK(clk), .Q(regs[42]) );
  DQV4_8TH40 regs_reg_30__9_ ( .D(n154), .CK(clk), .Q(regs[41]) );
  DQV4_8TH40 regs_reg_30__8_ ( .D(n153), .CK(clk), .Q(regs[40]) );
  DQV4_8TH40 regs_reg_30__7_ ( .D(n152), .CK(clk), .Q(regs[39]) );
  DQV4_8TH40 regs_reg_30__6_ ( .D(n151), .CK(clk), .Q(regs[38]) );
  DQV4_8TH40 regs_reg_30__5_ ( .D(n150), .CK(clk), .Q(regs[37]) );
  DQV4_8TH40 regs_reg_30__4_ ( .D(n149), .CK(clk), .Q(regs[36]) );
  DQV4_8TH40 regs_reg_30__3_ ( .D(n148), .CK(clk), .Q(regs[35]) );
  DQV4_8TH40 regs_reg_30__2_ ( .D(n147), .CK(clk), .Q(regs[34]) );
  DQV4_8TH40 regs_reg_30__1_ ( .D(n146), .CK(clk), .Q(regs[33]) );
  DQV4_8TH40 regs_reg_30__0_ ( .D(n145), .CK(clk), .Q(regs[32]) );
  DQV4_8TH40 regs_reg_31__31_ ( .D(n144), .CK(clk), .Q(regs[31]) );
  DQV4_8TH40 regs_reg_31__30_ ( .D(n143), .CK(clk), .Q(regs[30]) );
  DQV4_8TH40 regs_reg_31__29_ ( .D(n142), .CK(clk), .Q(regs[29]) );
  DQV4_8TH40 regs_reg_31__28_ ( .D(n141), .CK(clk), .Q(regs[28]) );
  DQV4_8TH40 regs_reg_31__27_ ( .D(n140), .CK(clk), .Q(regs[27]) );
  DQV4_8TH40 regs_reg_31__26_ ( .D(n139), .CK(clk), .Q(regs[26]) );
  DQV4_8TH40 regs_reg_31__25_ ( .D(n138), .CK(clk), .Q(regs[25]) );
  DQV4_8TH40 regs_reg_31__24_ ( .D(n137), .CK(clk), .Q(regs[24]) );
  DQV4_8TH40 regs_reg_31__23_ ( .D(n136), .CK(clk), .Q(regs[23]) );
  DQV4_8TH40 regs_reg_31__22_ ( .D(n135), .CK(clk), .Q(regs[22]) );
  DQV4_8TH40 regs_reg_31__21_ ( .D(n134), .CK(clk), .Q(regs[21]) );
  DQV4_8TH40 regs_reg_31__20_ ( .D(n133), .CK(clk), .Q(regs[20]) );
  DQV4_8TH40 regs_reg_31__19_ ( .D(n132), .CK(clk), .Q(regs[19]) );
  DQV4_8TH40 regs_reg_31__18_ ( .D(n131), .CK(clk), .Q(regs[18]) );
  DQV4_8TH40 regs_reg_31__17_ ( .D(n130), .CK(clk), .Q(regs[17]) );
  DQV4_8TH40 regs_reg_31__16_ ( .D(n129), .CK(clk), .Q(regs[16]) );
  DQV4_8TH40 regs_reg_31__15_ ( .D(n128), .CK(clk), .Q(regs[15]) );
  DQV4_8TH40 regs_reg_31__14_ ( .D(n127), .CK(clk), .Q(regs[14]) );
  DQV4_8TH40 regs_reg_31__13_ ( .D(n126), .CK(clk), .Q(regs[13]) );
  DQV4_8TH40 regs_reg_31__12_ ( .D(n125), .CK(clk), .Q(regs[12]) );
  DQV4_8TH40 regs_reg_31__11_ ( .D(n124), .CK(clk), .Q(regs[11]) );
  DQV4_8TH40 regs_reg_31__10_ ( .D(n123), .CK(clk), .Q(regs[10]) );
  DQV4_8TH40 regs_reg_31__9_ ( .D(n122), .CK(clk), .Q(regs[9]) );
  DQV4_8TH40 regs_reg_31__8_ ( .D(n121), .CK(clk), .Q(regs[8]) );
  DQV4_8TH40 regs_reg_31__7_ ( .D(n120), .CK(clk), .Q(regs[7]) );
  DQV4_8TH40 regs_reg_31__6_ ( .D(n119), .CK(clk), .Q(regs[6]) );
  DQV4_8TH40 regs_reg_31__5_ ( .D(n118), .CK(clk), .Q(regs[5]) );
  DQV4_8TH40 regs_reg_31__4_ ( .D(n117), .CK(clk), .Q(regs[4]) );
  DQV4_8TH40 regs_reg_31__3_ ( .D(n116), .CK(clk), .Q(regs[3]) );
  DQV4_8TH40 regs_reg_31__2_ ( .D(n115), .CK(clk), .Q(regs[2]) );
  DQV4_8TH40 regs_reg_31__1_ ( .D(n114), .CK(clk), .Q(regs[1]) );
  DQV4_8TH40 regs_reg_31__0_ ( .D(n113), .CK(clk), .Q(regs[0]) );
  EDQV2_8TH40 regs_reg_19__31_ ( .D(wdata[31]), .E(n1243), .CK(clk), .Q(
        regs[415]) );
  EDQV2_8TH40 regs_reg_19__30_ ( .D(wdata[30]), .E(n1243), .CK(clk), .Q(
        regs[414]) );
  EDQV2_8TH40 regs_reg_19__29_ ( .D(wdata[29]), .E(n1243), .CK(clk), .Q(
        regs[413]) );
  EDQV2_8TH40 regs_reg_19__28_ ( .D(wdata[28]), .E(n1243), .CK(clk), .Q(
        regs[412]) );
  EDQV2_8TH40 regs_reg_19__27_ ( .D(wdata[27]), .E(n1243), .CK(clk), .Q(
        regs[411]) );
  EDQV2_8TH40 regs_reg_19__26_ ( .D(wdata[26]), .E(n1243), .CK(clk), .Q(
        regs[410]) );
  EDQV2_8TH40 regs_reg_19__25_ ( .D(wdata[25]), .E(n1243), .CK(clk), .Q(
        regs[409]) );
  EDQV2_8TH40 regs_reg_19__24_ ( .D(wdata[24]), .E(n1243), .CK(clk), .Q(
        regs[408]) );
  EDQV2_8TH40 regs_reg_19__23_ ( .D(wdata[23]), .E(n1243), .CK(clk), .Q(
        regs[407]) );
  EDQV2_8TH40 regs_reg_19__22_ ( .D(wdata[22]), .E(n1243), .CK(clk), .Q(
        regs[406]) );
  EDQV2_8TH40 regs_reg_19__21_ ( .D(wdata[21]), .E(n1243), .CK(clk), .Q(
        regs[405]) );
  EDQV2_8TH40 regs_reg_19__20_ ( .D(wdata[20]), .E(n1243), .CK(clk), .Q(
        regs[404]) );
  EDQV2_8TH40 regs_reg_19__19_ ( .D(wdata[19]), .E(n1243), .CK(clk), .Q(
        regs[403]) );
  EDQV2_8TH40 regs_reg_19__18_ ( .D(wdata[18]), .E(n1243), .CK(clk), .Q(
        regs[402]) );
  EDQV2_8TH40 regs_reg_19__17_ ( .D(wdata[17]), .E(n1243), .CK(clk), .Q(
        regs[401]) );
  EDQV2_8TH40 regs_reg_19__16_ ( .D(wdata[16]), .E(n1243), .CK(clk), .Q(
        regs[400]) );
  EDQV2_8TH40 regs_reg_19__15_ ( .D(wdata[15]), .E(n1243), .CK(clk), .Q(
        regs[399]) );
  EDQV2_8TH40 regs_reg_19__14_ ( .D(wdata[14]), .E(n1243), .CK(clk), .Q(
        regs[398]) );
  EDQV2_8TH40 regs_reg_19__13_ ( .D(wdata[13]), .E(n1243), .CK(clk), .Q(
        regs[397]) );
  EDQV2_8TH40 regs_reg_19__12_ ( .D(wdata[12]), .E(n1243), .CK(clk), .Q(
        regs[396]) );
  EDQV2_8TH40 regs_reg_19__11_ ( .D(wdata[11]), .E(n1243), .CK(clk), .Q(
        regs[395]) );
  EDQV2_8TH40 regs_reg_19__10_ ( .D(wdata[10]), .E(n1243), .CK(clk), .Q(
        regs[394]) );
  EDQV2_8TH40 regs_reg_19__9_ ( .D(wdata[9]), .E(n1243), .CK(clk), .Q(
        regs[393]) );
  EDQV2_8TH40 regs_reg_19__8_ ( .D(wdata[8]), .E(n1243), .CK(clk), .Q(
        regs[392]) );
  EDQV2_8TH40 regs_reg_19__7_ ( .D(wdata[7]), .E(n1243), .CK(clk), .Q(
        regs[391]) );
  EDQV2_8TH40 regs_reg_19__6_ ( .D(wdata[6]), .E(n1243), .CK(clk), .Q(
        regs[390]) );
  EDQV2_8TH40 regs_reg_19__5_ ( .D(wdata[5]), .E(n1243), .CK(clk), .Q(
        regs[389]) );
  EDQV2_8TH40 regs_reg_19__4_ ( .D(wdata[4]), .E(n1243), .CK(clk), .Q(
        regs[388]) );
  EDQV2_8TH40 regs_reg_19__3_ ( .D(wdata[3]), .E(n1243), .CK(clk), .Q(
        regs[387]) );
  EDQV2_8TH40 regs_reg_19__2_ ( .D(wdata[2]), .E(n1243), .CK(clk), .Q(
        regs[386]) );
  EDQV2_8TH40 regs_reg_19__1_ ( .D(wdata[1]), .E(n1243), .CK(clk), .Q(
        regs[385]) );
  EDQV2_8TH40 regs_reg_19__0_ ( .D(wdata[0]), .E(n1243), .CK(clk), .Q(
        regs[384]) );
  EDQV2_8TH40 regs_reg_2__31_ ( .D(wdata[31]), .E(n1234), .CK(clk), .Q(
        regs[959]) );
  EDQV2_8TH40 regs_reg_2__30_ ( .D(wdata[30]), .E(n1234), .CK(clk), .Q(
        regs[958]) );
  EDQV2_8TH40 regs_reg_2__29_ ( .D(wdata[29]), .E(n1234), .CK(clk), .Q(
        regs[957]) );
  EDQV2_8TH40 regs_reg_2__28_ ( .D(wdata[28]), .E(n1234), .CK(clk), .Q(
        regs[956]) );
  EDQV2_8TH40 regs_reg_2__27_ ( .D(wdata[27]), .E(n1234), .CK(clk), .Q(
        regs[955]) );
  EDQV2_8TH40 regs_reg_2__26_ ( .D(wdata[26]), .E(n1234), .CK(clk), .Q(
        regs[954]) );
  EDQV2_8TH40 regs_reg_2__25_ ( .D(wdata[25]), .E(n1234), .CK(clk), .Q(
        regs[953]) );
  EDQV2_8TH40 regs_reg_2__24_ ( .D(wdata[24]), .E(n1234), .CK(clk), .Q(
        regs[952]) );
  EDQV2_8TH40 regs_reg_2__23_ ( .D(wdata[23]), .E(n1234), .CK(clk), .Q(
        regs[951]) );
  EDQV2_8TH40 regs_reg_2__22_ ( .D(wdata[22]), .E(n1234), .CK(clk), .Q(
        regs[950]) );
  EDQV2_8TH40 regs_reg_2__21_ ( .D(wdata[21]), .E(n1234), .CK(clk), .Q(
        regs[949]) );
  EDQV2_8TH40 regs_reg_2__20_ ( .D(wdata[20]), .E(n1234), .CK(clk), .Q(
        regs[948]) );
  EDQV2_8TH40 regs_reg_2__19_ ( .D(wdata[19]), .E(n1234), .CK(clk), .Q(
        regs[947]) );
  EDQV2_8TH40 regs_reg_2__18_ ( .D(wdata[18]), .E(n1234), .CK(clk), .Q(
        regs[946]) );
  EDQV2_8TH40 regs_reg_2__17_ ( .D(wdata[17]), .E(n1234), .CK(clk), .Q(
        regs[945]) );
  EDQV2_8TH40 regs_reg_2__16_ ( .D(wdata[16]), .E(n1234), .CK(clk), .Q(
        regs[944]) );
  EDQV2_8TH40 regs_reg_2__15_ ( .D(wdata[15]), .E(n1234), .CK(clk), .Q(
        regs[943]) );
  EDQV2_8TH40 regs_reg_2__14_ ( .D(wdata[14]), .E(n1234), .CK(clk), .Q(
        regs[942]) );
  EDQV2_8TH40 regs_reg_2__13_ ( .D(wdata[13]), .E(n1234), .CK(clk), .Q(
        regs[941]) );
  EDQV2_8TH40 regs_reg_2__12_ ( .D(wdata[12]), .E(n1234), .CK(clk), .Q(
        regs[940]) );
  EDQV2_8TH40 regs_reg_2__11_ ( .D(wdata[11]), .E(n1234), .CK(clk), .Q(
        regs[939]) );
  EDQV2_8TH40 regs_reg_2__10_ ( .D(wdata[10]), .E(n1234), .CK(clk), .Q(
        regs[938]) );
  EDQV2_8TH40 regs_reg_2__9_ ( .D(wdata[9]), .E(n1234), .CK(clk), .Q(regs[937]) );
  EDQV2_8TH40 regs_reg_2__8_ ( .D(wdata[8]), .E(n1234), .CK(clk), .Q(regs[936]) );
  EDQV2_8TH40 regs_reg_2__7_ ( .D(wdata[7]), .E(n1234), .CK(clk), .Q(regs[935]) );
  EDQV2_8TH40 regs_reg_2__6_ ( .D(wdata[6]), .E(n1234), .CK(clk), .Q(regs[934]) );
  EDQV2_8TH40 regs_reg_2__5_ ( .D(wdata[5]), .E(n1234), .CK(clk), .Q(regs[933]) );
  EDQV2_8TH40 regs_reg_2__4_ ( .D(wdata[4]), .E(n1234), .CK(clk), .Q(regs[932]) );
  EDQV2_8TH40 regs_reg_2__3_ ( .D(wdata[3]), .E(n1234), .CK(clk), .Q(regs[931]) );
  EDQV2_8TH40 regs_reg_2__2_ ( .D(wdata[2]), .E(n1234), .CK(clk), .Q(regs[930]) );
  EDQV2_8TH40 regs_reg_2__1_ ( .D(wdata[1]), .E(n1234), .CK(clk), .Q(regs[929]) );
  EDQV2_8TH40 regs_reg_2__0_ ( .D(wdata[0]), .E(n1234), .CK(clk), .Q(regs[928]) );
  EDQV2_8TH40 regs_reg_10__31_ ( .D(wdata[31]), .E(n1238), .CK(clk), .Q(
        regs[703]) );
  EDQV2_8TH40 regs_reg_10__30_ ( .D(wdata[30]), .E(n1238), .CK(clk), .Q(
        regs[702]) );
  EDQV2_8TH40 regs_reg_10__29_ ( .D(wdata[29]), .E(n1238), .CK(clk), .Q(
        regs[701]) );
  EDQV2_8TH40 regs_reg_10__28_ ( .D(wdata[28]), .E(n1238), .CK(clk), .Q(
        regs[700]) );
  EDQV2_8TH40 regs_reg_10__27_ ( .D(wdata[27]), .E(n1238), .CK(clk), .Q(
        regs[699]) );
  EDQV2_8TH40 regs_reg_10__26_ ( .D(wdata[26]), .E(n1238), .CK(clk), .Q(
        regs[698]) );
  EDQV2_8TH40 regs_reg_10__25_ ( .D(wdata[25]), .E(n1238), .CK(clk), .Q(
        regs[697]) );
  EDQV2_8TH40 regs_reg_10__24_ ( .D(wdata[24]), .E(n1238), .CK(clk), .Q(
        regs[696]) );
  EDQV2_8TH40 regs_reg_10__23_ ( .D(wdata[23]), .E(n1238), .CK(clk), .Q(
        regs[695]) );
  EDQV2_8TH40 regs_reg_10__22_ ( .D(wdata[22]), .E(n1238), .CK(clk), .Q(
        regs[694]) );
  EDQV2_8TH40 regs_reg_10__21_ ( .D(wdata[21]), .E(n1238), .CK(clk), .Q(
        regs[693]) );
  EDQV2_8TH40 regs_reg_10__20_ ( .D(wdata[20]), .E(n1238), .CK(clk), .Q(
        regs[692]) );
  EDQV2_8TH40 regs_reg_10__19_ ( .D(wdata[19]), .E(n1238), .CK(clk), .Q(
        regs[691]) );
  EDQV2_8TH40 regs_reg_10__18_ ( .D(wdata[18]), .E(n1238), .CK(clk), .Q(
        regs[690]) );
  EDQV2_8TH40 regs_reg_10__17_ ( .D(wdata[17]), .E(n1238), .CK(clk), .Q(
        regs[689]) );
  EDQV2_8TH40 regs_reg_10__16_ ( .D(wdata[16]), .E(n1238), .CK(clk), .Q(
        regs[688]) );
  EDQV2_8TH40 regs_reg_10__15_ ( .D(wdata[15]), .E(n1238), .CK(clk), .Q(
        regs[687]) );
  EDQV2_8TH40 regs_reg_10__14_ ( .D(wdata[14]), .E(n1238), .CK(clk), .Q(
        regs[686]) );
  EDQV2_8TH40 regs_reg_10__13_ ( .D(wdata[13]), .E(n1238), .CK(clk), .Q(
        regs[685]) );
  EDQV2_8TH40 regs_reg_10__12_ ( .D(wdata[12]), .E(n1238), .CK(clk), .Q(
        regs[684]) );
  EDQV2_8TH40 regs_reg_10__11_ ( .D(wdata[11]), .E(n1238), .CK(clk), .Q(
        regs[683]) );
  EDQV2_8TH40 regs_reg_10__10_ ( .D(wdata[10]), .E(n1238), .CK(clk), .Q(
        regs[682]) );
  EDQV2_8TH40 regs_reg_10__9_ ( .D(wdata[9]), .E(n1238), .CK(clk), .Q(
        regs[681]) );
  EDQV2_8TH40 regs_reg_10__8_ ( .D(wdata[8]), .E(n1238), .CK(clk), .Q(
        regs[680]) );
  EDQV2_8TH40 regs_reg_10__7_ ( .D(wdata[7]), .E(n1238), .CK(clk), .Q(
        regs[679]) );
  EDQV2_8TH40 regs_reg_10__6_ ( .D(wdata[6]), .E(n1238), .CK(clk), .Q(
        regs[678]) );
  EDQV2_8TH40 regs_reg_10__5_ ( .D(wdata[5]), .E(n1238), .CK(clk), .Q(
        regs[677]) );
  EDQV2_8TH40 regs_reg_10__4_ ( .D(wdata[4]), .E(n1238), .CK(clk), .Q(
        regs[676]) );
  EDQV2_8TH40 regs_reg_10__3_ ( .D(wdata[3]), .E(n1238), .CK(clk), .Q(
        regs[675]) );
  EDQV2_8TH40 regs_reg_10__2_ ( .D(wdata[2]), .E(n1238), .CK(clk), .Q(
        regs[674]) );
  EDQV2_8TH40 regs_reg_10__1_ ( .D(wdata[1]), .E(n1238), .CK(clk), .Q(
        regs[673]) );
  EDQV2_8TH40 regs_reg_10__0_ ( .D(wdata[0]), .E(n1238), .CK(clk), .Q(
        regs[672]) );
  EDQV2_8TH40 regs_reg_18__31_ ( .D(wdata[31]), .E(n1242), .CK(clk), .Q(
        regs[447]) );
  EDQV2_8TH40 regs_reg_18__30_ ( .D(wdata[30]), .E(n1242), .CK(clk), .Q(
        regs[446]) );
  EDQV2_8TH40 regs_reg_18__29_ ( .D(wdata[29]), .E(n1242), .CK(clk), .Q(
        regs[445]) );
  EDQV2_8TH40 regs_reg_18__28_ ( .D(wdata[28]), .E(n1242), .CK(clk), .Q(
        regs[444]) );
  EDQV2_8TH40 regs_reg_18__27_ ( .D(wdata[27]), .E(n1242), .CK(clk), .Q(
        regs[443]) );
  EDQV2_8TH40 regs_reg_18__26_ ( .D(wdata[26]), .E(n1242), .CK(clk), .Q(
        regs[442]) );
  EDQV2_8TH40 regs_reg_18__25_ ( .D(wdata[25]), .E(n1242), .CK(clk), .Q(
        regs[441]) );
  EDQV2_8TH40 regs_reg_18__24_ ( .D(wdata[24]), .E(n1242), .CK(clk), .Q(
        regs[440]) );
  EDQV2_8TH40 regs_reg_18__23_ ( .D(wdata[23]), .E(n1242), .CK(clk), .Q(
        regs[439]) );
  EDQV2_8TH40 regs_reg_18__22_ ( .D(wdata[22]), .E(n1242), .CK(clk), .Q(
        regs[438]) );
  EDQV2_8TH40 regs_reg_18__21_ ( .D(wdata[21]), .E(n1242), .CK(clk), .Q(
        regs[437]) );
  EDQV2_8TH40 regs_reg_18__20_ ( .D(wdata[20]), .E(n1242), .CK(clk), .Q(
        regs[436]) );
  EDQV2_8TH40 regs_reg_18__19_ ( .D(wdata[19]), .E(n1242), .CK(clk), .Q(
        regs[435]) );
  EDQV2_8TH40 regs_reg_18__18_ ( .D(wdata[18]), .E(n1242), .CK(clk), .Q(
        regs[434]) );
  EDQV2_8TH40 regs_reg_18__17_ ( .D(wdata[17]), .E(n1242), .CK(clk), .Q(
        regs[433]) );
  EDQV2_8TH40 regs_reg_18__16_ ( .D(wdata[16]), .E(n1242), .CK(clk), .Q(
        regs[432]) );
  EDQV2_8TH40 regs_reg_18__15_ ( .D(wdata[15]), .E(n1242), .CK(clk), .Q(
        regs[431]) );
  EDQV2_8TH40 regs_reg_18__14_ ( .D(wdata[14]), .E(n1242), .CK(clk), .Q(
        regs[430]) );
  EDQV2_8TH40 regs_reg_18__13_ ( .D(wdata[13]), .E(n1242), .CK(clk), .Q(
        regs[429]) );
  EDQV2_8TH40 regs_reg_18__12_ ( .D(wdata[12]), .E(n1242), .CK(clk), .Q(
        regs[428]) );
  EDQV2_8TH40 regs_reg_18__11_ ( .D(wdata[11]), .E(n1242), .CK(clk), .Q(
        regs[427]) );
  EDQV2_8TH40 regs_reg_18__10_ ( .D(wdata[10]), .E(n1242), .CK(clk), .Q(
        regs[426]) );
  EDQV2_8TH40 regs_reg_18__9_ ( .D(wdata[9]), .E(n1242), .CK(clk), .Q(
        regs[425]) );
  EDQV2_8TH40 regs_reg_18__8_ ( .D(wdata[8]), .E(n1242), .CK(clk), .Q(
        regs[424]) );
  EDQV2_8TH40 regs_reg_18__7_ ( .D(wdata[7]), .E(n1242), .CK(clk), .Q(
        regs[423]) );
  EDQV2_8TH40 regs_reg_18__6_ ( .D(wdata[6]), .E(n1242), .CK(clk), .Q(
        regs[422]) );
  EDQV2_8TH40 regs_reg_18__5_ ( .D(wdata[5]), .E(n1242), .CK(clk), .Q(
        regs[421]) );
  EDQV2_8TH40 regs_reg_18__4_ ( .D(wdata[4]), .E(n1242), .CK(clk), .Q(
        regs[420]) );
  EDQV2_8TH40 regs_reg_18__3_ ( .D(wdata[3]), .E(n1242), .CK(clk), .Q(
        regs[419]) );
  EDQV2_8TH40 regs_reg_18__2_ ( .D(wdata[2]), .E(n1242), .CK(clk), .Q(
        regs[418]) );
  EDQV2_8TH40 regs_reg_18__1_ ( .D(wdata[1]), .E(n1242), .CK(clk), .Q(
        regs[417]) );
  EDQV2_8TH40 regs_reg_18__0_ ( .D(wdata[0]), .E(n1242), .CK(clk), .Q(
        regs[416]) );
  EDQV2_8TH40 regs_reg_22__31_ ( .D(wdata[31]), .E(n1246), .CK(clk), .Q(
        regs[319]) );
  EDQV2_8TH40 regs_reg_22__30_ ( .D(wdata[30]), .E(n1246), .CK(clk), .Q(
        regs[318]) );
  EDQV2_8TH40 regs_reg_22__29_ ( .D(wdata[29]), .E(n1246), .CK(clk), .Q(
        regs[317]) );
  EDQV2_8TH40 regs_reg_22__28_ ( .D(wdata[28]), .E(n1246), .CK(clk), .Q(
        regs[316]) );
  EDQV2_8TH40 regs_reg_22__27_ ( .D(wdata[27]), .E(n1246), .CK(clk), .Q(
        regs[315]) );
  EDQV2_8TH40 regs_reg_22__26_ ( .D(wdata[26]), .E(n1246), .CK(clk), .Q(
        regs[314]) );
  EDQV2_8TH40 regs_reg_22__25_ ( .D(wdata[25]), .E(n1246), .CK(clk), .Q(
        regs[313]) );
  EDQV2_8TH40 regs_reg_22__24_ ( .D(wdata[24]), .E(n1246), .CK(clk), .Q(
        regs[312]) );
  EDQV2_8TH40 regs_reg_22__23_ ( .D(wdata[23]), .E(n1246), .CK(clk), .Q(
        regs[311]) );
  EDQV2_8TH40 regs_reg_22__22_ ( .D(wdata[22]), .E(n1246), .CK(clk), .Q(
        regs[310]) );
  EDQV2_8TH40 regs_reg_22__21_ ( .D(wdata[21]), .E(n1246), .CK(clk), .Q(
        regs[309]) );
  EDQV2_8TH40 regs_reg_22__20_ ( .D(wdata[20]), .E(n1246), .CK(clk), .Q(
        regs[308]) );
  EDQV2_8TH40 regs_reg_22__19_ ( .D(wdata[19]), .E(n1246), .CK(clk), .Q(
        regs[307]) );
  EDQV2_8TH40 regs_reg_22__18_ ( .D(wdata[18]), .E(n1246), .CK(clk), .Q(
        regs[306]) );
  EDQV2_8TH40 regs_reg_22__17_ ( .D(wdata[17]), .E(n1246), .CK(clk), .Q(
        regs[305]) );
  EDQV2_8TH40 regs_reg_22__16_ ( .D(wdata[16]), .E(n1246), .CK(clk), .Q(
        regs[304]) );
  EDQV2_8TH40 regs_reg_22__15_ ( .D(wdata[15]), .E(n1246), .CK(clk), .Q(
        regs[303]) );
  EDQV2_8TH40 regs_reg_22__14_ ( .D(wdata[14]), .E(n1246), .CK(clk), .Q(
        regs[302]) );
  EDQV2_8TH40 regs_reg_22__13_ ( .D(wdata[13]), .E(n1246), .CK(clk), .Q(
        regs[301]) );
  EDQV2_8TH40 regs_reg_22__12_ ( .D(wdata[12]), .E(n1246), .CK(clk), .Q(
        regs[300]) );
  EDQV2_8TH40 regs_reg_22__11_ ( .D(wdata[11]), .E(n1246), .CK(clk), .Q(
        regs[299]) );
  EDQV2_8TH40 regs_reg_22__10_ ( .D(wdata[10]), .E(n1246), .CK(clk), .Q(
        regs[298]) );
  EDQV2_8TH40 regs_reg_22__9_ ( .D(wdata[9]), .E(n1246), .CK(clk), .Q(
        regs[297]) );
  EDQV2_8TH40 regs_reg_22__8_ ( .D(wdata[8]), .E(n1246), .CK(clk), .Q(
        regs[296]) );
  EDQV2_8TH40 regs_reg_22__7_ ( .D(wdata[7]), .E(n1246), .CK(clk), .Q(
        regs[295]) );
  EDQV2_8TH40 regs_reg_22__6_ ( .D(wdata[6]), .E(n1246), .CK(clk), .Q(
        regs[294]) );
  EDQV2_8TH40 regs_reg_22__5_ ( .D(wdata[5]), .E(n1246), .CK(clk), .Q(
        regs[293]) );
  EDQV2_8TH40 regs_reg_22__4_ ( .D(wdata[4]), .E(n1246), .CK(clk), .Q(
        regs[292]) );
  EDQV2_8TH40 regs_reg_22__3_ ( .D(wdata[3]), .E(n1246), .CK(clk), .Q(
        regs[291]) );
  EDQV2_8TH40 regs_reg_22__2_ ( .D(wdata[2]), .E(n1246), .CK(clk), .Q(
        regs[290]) );
  EDQV2_8TH40 regs_reg_22__1_ ( .D(wdata[1]), .E(n1246), .CK(clk), .Q(
        regs[289]) );
  EDQV2_8TH40 regs_reg_22__0_ ( .D(wdata[0]), .E(n1246), .CK(clk), .Q(
        regs[288]) );
  EDQV2_8TH40 regs_reg_26__31_ ( .D(wdata[31]), .E(n1249), .CK(clk), .Q(
        regs[191]) );
  EDQV2_8TH40 regs_reg_26__30_ ( .D(wdata[30]), .E(n1249), .CK(clk), .Q(
        regs[190]) );
  EDQV2_8TH40 regs_reg_26__29_ ( .D(wdata[29]), .E(n1249), .CK(clk), .Q(
        regs[189]) );
  EDQV2_8TH40 regs_reg_26__28_ ( .D(wdata[28]), .E(n1249), .CK(clk), .Q(
        regs[188]) );
  EDQV2_8TH40 regs_reg_26__27_ ( .D(wdata[27]), .E(n1249), .CK(clk), .Q(
        regs[187]) );
  EDQV2_8TH40 regs_reg_26__26_ ( .D(wdata[26]), .E(n1249), .CK(clk), .Q(
        regs[186]) );
  EDQV2_8TH40 regs_reg_26__25_ ( .D(wdata[25]), .E(n1249), .CK(clk), .Q(
        regs[185]) );
  EDQV2_8TH40 regs_reg_26__24_ ( .D(wdata[24]), .E(n1249), .CK(clk), .Q(
        regs[184]) );
  EDQV2_8TH40 regs_reg_26__23_ ( .D(wdata[23]), .E(n1249), .CK(clk), .Q(
        regs[183]) );
  EDQV2_8TH40 regs_reg_26__22_ ( .D(wdata[22]), .E(n1249), .CK(clk), .Q(
        regs[182]) );
  EDQV2_8TH40 regs_reg_26__21_ ( .D(wdata[21]), .E(n1249), .CK(clk), .Q(
        regs[181]) );
  EDQV2_8TH40 regs_reg_26__20_ ( .D(wdata[20]), .E(n1249), .CK(clk), .Q(
        regs[180]) );
  EDQV2_8TH40 regs_reg_26__19_ ( .D(wdata[19]), .E(n1249), .CK(clk), .Q(
        regs[179]) );
  EDQV2_8TH40 regs_reg_26__18_ ( .D(wdata[18]), .E(n1249), .CK(clk), .Q(
        regs[178]) );
  EDQV2_8TH40 regs_reg_26__17_ ( .D(wdata[17]), .E(n1249), .CK(clk), .Q(
        regs[177]) );
  EDQV2_8TH40 regs_reg_26__16_ ( .D(wdata[16]), .E(n1249), .CK(clk), .Q(
        regs[176]) );
  EDQV2_8TH40 regs_reg_26__15_ ( .D(wdata[15]), .E(n1249), .CK(clk), .Q(
        regs[175]) );
  EDQV2_8TH40 regs_reg_26__14_ ( .D(wdata[14]), .E(n1249), .CK(clk), .Q(
        regs[174]) );
  EDQV2_8TH40 regs_reg_26__13_ ( .D(wdata[13]), .E(n1249), .CK(clk), .Q(
        regs[173]) );
  EDQV2_8TH40 regs_reg_26__12_ ( .D(wdata[12]), .E(n1249), .CK(clk), .Q(
        regs[172]) );
  EDQV2_8TH40 regs_reg_26__11_ ( .D(wdata[11]), .E(n1249), .CK(clk), .Q(
        regs[171]) );
  EDQV2_8TH40 regs_reg_26__10_ ( .D(wdata[10]), .E(n1249), .CK(clk), .Q(
        regs[170]) );
  EDQV2_8TH40 regs_reg_26__9_ ( .D(wdata[9]), .E(n1249), .CK(clk), .Q(
        regs[169]) );
  EDQV2_8TH40 regs_reg_26__8_ ( .D(wdata[8]), .E(n1249), .CK(clk), .Q(
        regs[168]) );
  EDQV2_8TH40 regs_reg_26__7_ ( .D(wdata[7]), .E(n1249), .CK(clk), .Q(
        regs[167]) );
  EDQV2_8TH40 regs_reg_26__6_ ( .D(wdata[6]), .E(n1249), .CK(clk), .Q(
        regs[166]) );
  EDQV2_8TH40 regs_reg_26__5_ ( .D(wdata[5]), .E(n1249), .CK(clk), .Q(
        regs[165]) );
  EDQV2_8TH40 regs_reg_26__4_ ( .D(wdata[4]), .E(n1249), .CK(clk), .Q(
        regs[164]) );
  EDQV2_8TH40 regs_reg_26__3_ ( .D(wdata[3]), .E(n1249), .CK(clk), .Q(
        regs[163]) );
  EDQV2_8TH40 regs_reg_26__2_ ( .D(wdata[2]), .E(n1249), .CK(clk), .Q(
        regs[162]) );
  EDQV2_8TH40 regs_reg_26__1_ ( .D(wdata[1]), .E(n1249), .CK(clk), .Q(
        regs[161]) );
  EDQV2_8TH40 regs_reg_26__0_ ( .D(wdata[0]), .E(n1249), .CK(clk), .Q(
        regs[160]) );
  EDQV2_8TH40 regs_reg_4__31_ ( .D(wdata[31]), .E(n1235), .CK(clk), .Q(
        regs[895]) );
  EDQV2_8TH40 regs_reg_4__30_ ( .D(wdata[30]), .E(n1235), .CK(clk), .Q(
        regs[894]) );
  EDQV2_8TH40 regs_reg_4__29_ ( .D(wdata[29]), .E(n1235), .CK(clk), .Q(
        regs[893]) );
  EDQV2_8TH40 regs_reg_4__28_ ( .D(wdata[28]), .E(n1235), .CK(clk), .Q(
        regs[892]) );
  EDQV2_8TH40 regs_reg_4__27_ ( .D(wdata[27]), .E(n1235), .CK(clk), .Q(
        regs[891]) );
  EDQV2_8TH40 regs_reg_4__26_ ( .D(wdata[26]), .E(n1235), .CK(clk), .Q(
        regs[890]) );
  EDQV2_8TH40 regs_reg_4__25_ ( .D(wdata[25]), .E(n1235), .CK(clk), .Q(
        regs[889]) );
  EDQV2_8TH40 regs_reg_4__24_ ( .D(wdata[24]), .E(n1235), .CK(clk), .Q(
        regs[888]) );
  EDQV2_8TH40 regs_reg_4__23_ ( .D(wdata[23]), .E(n1235), .CK(clk), .Q(
        regs[887]) );
  EDQV2_8TH40 regs_reg_4__22_ ( .D(wdata[22]), .E(n1235), .CK(clk), .Q(
        regs[886]) );
  EDQV2_8TH40 regs_reg_4__21_ ( .D(wdata[21]), .E(n1235), .CK(clk), .Q(
        regs[885]) );
  EDQV2_8TH40 regs_reg_4__20_ ( .D(wdata[20]), .E(n1235), .CK(clk), .Q(
        regs[884]) );
  EDQV2_8TH40 regs_reg_4__19_ ( .D(wdata[19]), .E(n1235), .CK(clk), .Q(
        regs[883]) );
  EDQV2_8TH40 regs_reg_4__18_ ( .D(wdata[18]), .E(n1235), .CK(clk), .Q(
        regs[882]) );
  EDQV2_8TH40 regs_reg_4__17_ ( .D(wdata[17]), .E(n1235), .CK(clk), .Q(
        regs[881]) );
  EDQV2_8TH40 regs_reg_4__16_ ( .D(wdata[16]), .E(n1235), .CK(clk), .Q(
        regs[880]) );
  EDQV2_8TH40 regs_reg_4__15_ ( .D(wdata[15]), .E(n1235), .CK(clk), .Q(
        regs[879]) );
  EDQV2_8TH40 regs_reg_4__14_ ( .D(wdata[14]), .E(n1235), .CK(clk), .Q(
        regs[878]) );
  EDQV2_8TH40 regs_reg_4__13_ ( .D(wdata[13]), .E(n1235), .CK(clk), .Q(
        regs[877]) );
  EDQV2_8TH40 regs_reg_4__12_ ( .D(wdata[12]), .E(n1235), .CK(clk), .Q(
        regs[876]) );
  EDQV2_8TH40 regs_reg_4__11_ ( .D(wdata[11]), .E(n1235), .CK(clk), .Q(
        regs[875]) );
  EDQV2_8TH40 regs_reg_4__10_ ( .D(wdata[10]), .E(n1235), .CK(clk), .Q(
        regs[874]) );
  EDQV2_8TH40 regs_reg_4__9_ ( .D(wdata[9]), .E(n1235), .CK(clk), .Q(regs[873]) );
  EDQV2_8TH40 regs_reg_4__8_ ( .D(wdata[8]), .E(n1235), .CK(clk), .Q(regs[872]) );
  EDQV2_8TH40 regs_reg_4__7_ ( .D(wdata[7]), .E(n1235), .CK(clk), .Q(regs[871]) );
  EDQV2_8TH40 regs_reg_4__6_ ( .D(wdata[6]), .E(n1235), .CK(clk), .Q(regs[870]) );
  EDQV2_8TH40 regs_reg_4__5_ ( .D(wdata[5]), .E(n1235), .CK(clk), .Q(regs[869]) );
  EDQV2_8TH40 regs_reg_4__4_ ( .D(wdata[4]), .E(n1235), .CK(clk), .Q(regs[868]) );
  EDQV2_8TH40 regs_reg_4__3_ ( .D(wdata[3]), .E(n1235), .CK(clk), .Q(regs[867]) );
  EDQV2_8TH40 regs_reg_4__2_ ( .D(wdata[2]), .E(n1235), .CK(clk), .Q(regs[866]) );
  EDQV2_8TH40 regs_reg_4__1_ ( .D(wdata[1]), .E(n1235), .CK(clk), .Q(regs[865]) );
  EDQV2_8TH40 regs_reg_4__0_ ( .D(wdata[0]), .E(n1235), .CK(clk), .Q(regs[864]) );
  EDQV2_8TH40 regs_reg_8__31_ ( .D(wdata[31]), .E(n1236), .CK(clk), .Q(
        regs[767]) );
  EDQV2_8TH40 regs_reg_8__30_ ( .D(wdata[30]), .E(n1236), .CK(clk), .Q(
        regs[766]) );
  EDQV2_8TH40 regs_reg_8__29_ ( .D(wdata[29]), .E(n1236), .CK(clk), .Q(
        regs[765]) );
  EDQV2_8TH40 regs_reg_8__28_ ( .D(wdata[28]), .E(n1236), .CK(clk), .Q(
        regs[764]) );
  EDQV2_8TH40 regs_reg_8__27_ ( .D(wdata[27]), .E(n1236), .CK(clk), .Q(
        regs[763]) );
  EDQV2_8TH40 regs_reg_8__26_ ( .D(wdata[26]), .E(n1236), .CK(clk), .Q(
        regs[762]) );
  EDQV2_8TH40 regs_reg_8__25_ ( .D(wdata[25]), .E(n1236), .CK(clk), .Q(
        regs[761]) );
  EDQV2_8TH40 regs_reg_8__24_ ( .D(wdata[24]), .E(n1236), .CK(clk), .Q(
        regs[760]) );
  EDQV2_8TH40 regs_reg_8__23_ ( .D(wdata[23]), .E(n1236), .CK(clk), .Q(
        regs[759]) );
  EDQV2_8TH40 regs_reg_8__22_ ( .D(wdata[22]), .E(n1236), .CK(clk), .Q(
        regs[758]) );
  EDQV2_8TH40 regs_reg_8__21_ ( .D(wdata[21]), .E(n1236), .CK(clk), .Q(
        regs[757]) );
  EDQV2_8TH40 regs_reg_8__20_ ( .D(wdata[20]), .E(n1236), .CK(clk), .Q(
        regs[756]) );
  EDQV2_8TH40 regs_reg_8__19_ ( .D(wdata[19]), .E(n1236), .CK(clk), .Q(
        regs[755]) );
  EDQV2_8TH40 regs_reg_8__18_ ( .D(wdata[18]), .E(n1236), .CK(clk), .Q(
        regs[754]) );
  EDQV2_8TH40 regs_reg_8__17_ ( .D(wdata[17]), .E(n1236), .CK(clk), .Q(
        regs[753]) );
  EDQV2_8TH40 regs_reg_8__16_ ( .D(wdata[16]), .E(n1236), .CK(clk), .Q(
        regs[752]) );
  EDQV2_8TH40 regs_reg_8__15_ ( .D(wdata[15]), .E(n1236), .CK(clk), .Q(
        regs[751]) );
  EDQV2_8TH40 regs_reg_8__14_ ( .D(wdata[14]), .E(n1236), .CK(clk), .Q(
        regs[750]) );
  EDQV2_8TH40 regs_reg_8__13_ ( .D(wdata[13]), .E(n1236), .CK(clk), .Q(
        regs[749]) );
  EDQV2_8TH40 regs_reg_8__12_ ( .D(wdata[12]), .E(n1236), .CK(clk), .Q(
        regs[748]) );
  EDQV2_8TH40 regs_reg_8__11_ ( .D(wdata[11]), .E(n1236), .CK(clk), .Q(
        regs[747]) );
  EDQV2_8TH40 regs_reg_8__10_ ( .D(wdata[10]), .E(n1236), .CK(clk), .Q(
        regs[746]) );
  EDQV2_8TH40 regs_reg_8__9_ ( .D(wdata[9]), .E(n1236), .CK(clk), .Q(regs[745]) );
  EDQV2_8TH40 regs_reg_8__8_ ( .D(wdata[8]), .E(n1236), .CK(clk), .Q(regs[744]) );
  EDQV2_8TH40 regs_reg_8__7_ ( .D(wdata[7]), .E(n1236), .CK(clk), .Q(regs[743]) );
  EDQV2_8TH40 regs_reg_8__6_ ( .D(wdata[6]), .E(n1236), .CK(clk), .Q(regs[742]) );
  EDQV2_8TH40 regs_reg_8__5_ ( .D(wdata[5]), .E(n1236), .CK(clk), .Q(regs[741]) );
  EDQV2_8TH40 regs_reg_8__4_ ( .D(wdata[4]), .E(n1236), .CK(clk), .Q(regs[740]) );
  EDQV2_8TH40 regs_reg_8__3_ ( .D(wdata[3]), .E(n1236), .CK(clk), .Q(regs[739]) );
  EDQV2_8TH40 regs_reg_8__2_ ( .D(wdata[2]), .E(n1236), .CK(clk), .Q(regs[738]) );
  EDQV2_8TH40 regs_reg_8__1_ ( .D(wdata[1]), .E(n1236), .CK(clk), .Q(regs[737]) );
  EDQV2_8TH40 regs_reg_8__0_ ( .D(wdata[0]), .E(n1236), .CK(clk), .Q(regs[736]) );
  EDQV2_8TH40 regs_reg_12__31_ ( .D(wdata[31]), .E(n1239), .CK(clk), .Q(
        regs[639]) );
  EDQV2_8TH40 regs_reg_12__30_ ( .D(wdata[30]), .E(n1239), .CK(clk), .Q(
        regs[638]) );
  EDQV2_8TH40 regs_reg_12__29_ ( .D(wdata[29]), .E(n1239), .CK(clk), .Q(
        regs[637]) );
  EDQV2_8TH40 regs_reg_12__28_ ( .D(wdata[28]), .E(n1239), .CK(clk), .Q(
        regs[636]) );
  EDQV2_8TH40 regs_reg_12__27_ ( .D(wdata[27]), .E(n1239), .CK(clk), .Q(
        regs[635]) );
  EDQV2_8TH40 regs_reg_12__26_ ( .D(wdata[26]), .E(n1239), .CK(clk), .Q(
        regs[634]) );
  EDQV2_8TH40 regs_reg_12__25_ ( .D(wdata[25]), .E(n1239), .CK(clk), .Q(
        regs[633]) );
  EDQV2_8TH40 regs_reg_12__24_ ( .D(wdata[24]), .E(n1239), .CK(clk), .Q(
        regs[632]) );
  EDQV2_8TH40 regs_reg_12__23_ ( .D(wdata[23]), .E(n1239), .CK(clk), .Q(
        regs[631]) );
  EDQV2_8TH40 regs_reg_12__22_ ( .D(wdata[22]), .E(n1239), .CK(clk), .Q(
        regs[630]) );
  EDQV2_8TH40 regs_reg_12__21_ ( .D(wdata[21]), .E(n1239), .CK(clk), .Q(
        regs[629]) );
  EDQV2_8TH40 regs_reg_12__20_ ( .D(wdata[20]), .E(n1239), .CK(clk), .Q(
        regs[628]) );
  EDQV2_8TH40 regs_reg_12__19_ ( .D(wdata[19]), .E(n1239), .CK(clk), .Q(
        regs[627]) );
  EDQV2_8TH40 regs_reg_12__18_ ( .D(wdata[18]), .E(n1239), .CK(clk), .Q(
        regs[626]) );
  EDQV2_8TH40 regs_reg_12__17_ ( .D(wdata[17]), .E(n1239), .CK(clk), .Q(
        regs[625]) );
  EDQV2_8TH40 regs_reg_12__16_ ( .D(wdata[16]), .E(n1239), .CK(clk), .Q(
        regs[624]) );
  EDQV2_8TH40 regs_reg_12__15_ ( .D(wdata[15]), .E(n1239), .CK(clk), .Q(
        regs[623]) );
  EDQV2_8TH40 regs_reg_12__14_ ( .D(wdata[14]), .E(n1239), .CK(clk), .Q(
        regs[622]) );
  EDQV2_8TH40 regs_reg_12__13_ ( .D(wdata[13]), .E(n1239), .CK(clk), .Q(
        regs[621]) );
  EDQV2_8TH40 regs_reg_12__12_ ( .D(wdata[12]), .E(n1239), .CK(clk), .Q(
        regs[620]) );
  EDQV2_8TH40 regs_reg_12__11_ ( .D(wdata[11]), .E(n1239), .CK(clk), .Q(
        regs[619]) );
  EDQV2_8TH40 regs_reg_12__10_ ( .D(wdata[10]), .E(n1239), .CK(clk), .Q(
        regs[618]) );
  EDQV2_8TH40 regs_reg_12__9_ ( .D(wdata[9]), .E(n1239), .CK(clk), .Q(
        regs[617]) );
  EDQV2_8TH40 regs_reg_12__8_ ( .D(wdata[8]), .E(n1239), .CK(clk), .Q(
        regs[616]) );
  EDQV2_8TH40 regs_reg_12__7_ ( .D(wdata[7]), .E(n1239), .CK(clk), .Q(
        regs[615]) );
  EDQV2_8TH40 regs_reg_12__6_ ( .D(wdata[6]), .E(n1239), .CK(clk), .Q(
        regs[614]) );
  EDQV2_8TH40 regs_reg_12__5_ ( .D(wdata[5]), .E(n1239), .CK(clk), .Q(
        regs[613]) );
  EDQV2_8TH40 regs_reg_12__4_ ( .D(wdata[4]), .E(n1239), .CK(clk), .Q(
        regs[612]) );
  EDQV2_8TH40 regs_reg_12__3_ ( .D(wdata[3]), .E(n1239), .CK(clk), .Q(
        regs[611]) );
  EDQV2_8TH40 regs_reg_12__2_ ( .D(wdata[2]), .E(n1239), .CK(clk), .Q(
        regs[610]) );
  EDQV2_8TH40 regs_reg_12__1_ ( .D(wdata[1]), .E(n1239), .CK(clk), .Q(
        regs[609]) );
  EDQV2_8TH40 regs_reg_12__0_ ( .D(wdata[0]), .E(n1239), .CK(clk), .Q(
        regs[608]) );
  EDQV2_8TH40 regs_reg_16__31_ ( .D(wdata[31]), .E(n1240), .CK(clk), .Q(
        regs[511]) );
  EDQV2_8TH40 regs_reg_16__30_ ( .D(wdata[30]), .E(n1240), .CK(clk), .Q(
        regs[510]) );
  EDQV2_8TH40 regs_reg_16__29_ ( .D(wdata[29]), .E(n1240), .CK(clk), .Q(
        regs[509]) );
  EDQV2_8TH40 regs_reg_16__28_ ( .D(wdata[28]), .E(n1240), .CK(clk), .Q(
        regs[508]) );
  EDQV2_8TH40 regs_reg_16__27_ ( .D(wdata[27]), .E(n1240), .CK(clk), .Q(
        regs[507]) );
  EDQV2_8TH40 regs_reg_16__26_ ( .D(wdata[26]), .E(n1240), .CK(clk), .Q(
        regs[506]) );
  EDQV2_8TH40 regs_reg_16__25_ ( .D(wdata[25]), .E(n1240), .CK(clk), .Q(
        regs[505]) );
  EDQV2_8TH40 regs_reg_16__24_ ( .D(wdata[24]), .E(n1240), .CK(clk), .Q(
        regs[504]) );
  EDQV2_8TH40 regs_reg_16__23_ ( .D(wdata[23]), .E(n1240), .CK(clk), .Q(
        regs[503]) );
  EDQV2_8TH40 regs_reg_16__22_ ( .D(wdata[22]), .E(n1240), .CK(clk), .Q(
        regs[502]) );
  EDQV2_8TH40 regs_reg_16__21_ ( .D(wdata[21]), .E(n1240), .CK(clk), .Q(
        regs[501]) );
  EDQV2_8TH40 regs_reg_16__20_ ( .D(wdata[20]), .E(n1240), .CK(clk), .Q(
        regs[500]) );
  EDQV2_8TH40 regs_reg_16__19_ ( .D(wdata[19]), .E(n1240), .CK(clk), .Q(
        regs[499]) );
  EDQV2_8TH40 regs_reg_16__18_ ( .D(wdata[18]), .E(n1240), .CK(clk), .Q(
        regs[498]) );
  EDQV2_8TH40 regs_reg_16__17_ ( .D(wdata[17]), .E(n1240), .CK(clk), .Q(
        regs[497]) );
  EDQV2_8TH40 regs_reg_16__16_ ( .D(wdata[16]), .E(n1240), .CK(clk), .Q(
        regs[496]) );
  EDQV2_8TH40 regs_reg_16__15_ ( .D(wdata[15]), .E(n1240), .CK(clk), .Q(
        regs[495]) );
  EDQV2_8TH40 regs_reg_16__14_ ( .D(wdata[14]), .E(n1240), .CK(clk), .Q(
        regs[494]) );
  EDQV2_8TH40 regs_reg_16__13_ ( .D(wdata[13]), .E(n1240), .CK(clk), .Q(
        regs[493]) );
  EDQV2_8TH40 regs_reg_16__12_ ( .D(wdata[12]), .E(n1240), .CK(clk), .Q(
        regs[492]) );
  EDQV2_8TH40 regs_reg_16__11_ ( .D(wdata[11]), .E(n1240), .CK(clk), .Q(
        regs[491]) );
  EDQV2_8TH40 regs_reg_16__10_ ( .D(wdata[10]), .E(n1240), .CK(clk), .Q(
        regs[490]) );
  EDQV2_8TH40 regs_reg_16__9_ ( .D(wdata[9]), .E(n1240), .CK(clk), .Q(
        regs[489]) );
  EDQV2_8TH40 regs_reg_16__8_ ( .D(wdata[8]), .E(n1240), .CK(clk), .Q(
        regs[488]) );
  EDQV2_8TH40 regs_reg_16__7_ ( .D(wdata[7]), .E(n1240), .CK(clk), .Q(
        regs[487]) );
  EDQV2_8TH40 regs_reg_16__6_ ( .D(wdata[6]), .E(n1240), .CK(clk), .Q(
        regs[486]) );
  EDQV2_8TH40 regs_reg_16__5_ ( .D(wdata[5]), .E(n1240), .CK(clk), .Q(
        regs[485]) );
  EDQV2_8TH40 regs_reg_16__4_ ( .D(wdata[4]), .E(n1240), .CK(clk), .Q(
        regs[484]) );
  EDQV2_8TH40 regs_reg_16__3_ ( .D(wdata[3]), .E(n1240), .CK(clk), .Q(
        regs[483]) );
  EDQV2_8TH40 regs_reg_16__2_ ( .D(wdata[2]), .E(n1240), .CK(clk), .Q(
        regs[482]) );
  EDQV2_8TH40 regs_reg_16__1_ ( .D(wdata[1]), .E(n1240), .CK(clk), .Q(
        regs[481]) );
  EDQV2_8TH40 regs_reg_16__0_ ( .D(wdata[0]), .E(n1240), .CK(clk), .Q(
        regs[480]) );
  EDQV2_8TH40 regs_reg_20__31_ ( .D(wdata[31]), .E(n1244), .CK(clk), .Q(
        regs[383]) );
  EDQV2_8TH40 regs_reg_20__30_ ( .D(wdata[30]), .E(n1244), .CK(clk), .Q(
        regs[382]) );
  EDQV2_8TH40 regs_reg_20__29_ ( .D(wdata[29]), .E(n1244), .CK(clk), .Q(
        regs[381]) );
  EDQV2_8TH40 regs_reg_20__28_ ( .D(wdata[28]), .E(n1244), .CK(clk), .Q(
        regs[380]) );
  EDQV2_8TH40 regs_reg_20__27_ ( .D(wdata[27]), .E(n1244), .CK(clk), .Q(
        regs[379]) );
  EDQV2_8TH40 regs_reg_20__26_ ( .D(wdata[26]), .E(n1244), .CK(clk), .Q(
        regs[378]) );
  EDQV2_8TH40 regs_reg_20__25_ ( .D(wdata[25]), .E(n1244), .CK(clk), .Q(
        regs[377]) );
  EDQV2_8TH40 regs_reg_20__24_ ( .D(wdata[24]), .E(n1244), .CK(clk), .Q(
        regs[376]) );
  EDQV2_8TH40 regs_reg_20__23_ ( .D(wdata[23]), .E(n1244), .CK(clk), .Q(
        regs[375]) );
  EDQV2_8TH40 regs_reg_20__22_ ( .D(wdata[22]), .E(n1244), .CK(clk), .Q(
        regs[374]) );
  EDQV2_8TH40 regs_reg_20__21_ ( .D(wdata[21]), .E(n1244), .CK(clk), .Q(
        regs[373]) );
  EDQV2_8TH40 regs_reg_20__20_ ( .D(wdata[20]), .E(n1244), .CK(clk), .Q(
        regs[372]) );
  EDQV2_8TH40 regs_reg_20__19_ ( .D(wdata[19]), .E(n1244), .CK(clk), .Q(
        regs[371]) );
  EDQV2_8TH40 regs_reg_20__18_ ( .D(wdata[18]), .E(n1244), .CK(clk), .Q(
        regs[370]) );
  EDQV2_8TH40 regs_reg_20__17_ ( .D(wdata[17]), .E(n1244), .CK(clk), .Q(
        regs[369]) );
  EDQV2_8TH40 regs_reg_20__16_ ( .D(wdata[16]), .E(n1244), .CK(clk), .Q(
        regs[368]) );
  EDQV2_8TH40 regs_reg_20__15_ ( .D(wdata[15]), .E(n1244), .CK(clk), .Q(
        regs[367]) );
  EDQV2_8TH40 regs_reg_20__14_ ( .D(wdata[14]), .E(n1244), .CK(clk), .Q(
        regs[366]) );
  EDQV2_8TH40 regs_reg_20__13_ ( .D(wdata[13]), .E(n1244), .CK(clk), .Q(
        regs[365]) );
  EDQV2_8TH40 regs_reg_20__12_ ( .D(wdata[12]), .E(n1244), .CK(clk), .Q(
        regs[364]) );
  EDQV2_8TH40 regs_reg_20__11_ ( .D(wdata[11]), .E(n1244), .CK(clk), .Q(
        regs[363]) );
  EDQV2_8TH40 regs_reg_20__10_ ( .D(wdata[10]), .E(n1244), .CK(clk), .Q(
        regs[362]) );
  EDQV2_8TH40 regs_reg_20__9_ ( .D(wdata[9]), .E(n1244), .CK(clk), .Q(
        regs[361]) );
  EDQV2_8TH40 regs_reg_20__8_ ( .D(wdata[8]), .E(n1244), .CK(clk), .Q(
        regs[360]) );
  EDQV2_8TH40 regs_reg_20__7_ ( .D(wdata[7]), .E(n1244), .CK(clk), .Q(
        regs[359]) );
  EDQV2_8TH40 regs_reg_20__6_ ( .D(wdata[6]), .E(n1244), .CK(clk), .Q(
        regs[358]) );
  EDQV2_8TH40 regs_reg_20__5_ ( .D(wdata[5]), .E(n1244), .CK(clk), .Q(
        regs[357]) );
  EDQV2_8TH40 regs_reg_20__4_ ( .D(wdata[4]), .E(n1244), .CK(clk), .Q(
        regs[356]) );
  EDQV2_8TH40 regs_reg_20__3_ ( .D(wdata[3]), .E(n1244), .CK(clk), .Q(
        regs[355]) );
  EDQV2_8TH40 regs_reg_20__2_ ( .D(wdata[2]), .E(n1244), .CK(clk), .Q(
        regs[354]) );
  EDQV2_8TH40 regs_reg_20__1_ ( .D(wdata[1]), .E(n1244), .CK(clk), .Q(
        regs[353]) );
  EDQV2_8TH40 regs_reg_20__0_ ( .D(wdata[0]), .E(n1244), .CK(clk), .Q(
        regs[352]) );
  EDQV2_8TH40 regs_reg_24__31_ ( .D(wdata[31]), .E(n1247), .CK(clk), .Q(
        regs[255]) );
  EDQV2_8TH40 regs_reg_24__30_ ( .D(wdata[30]), .E(n1247), .CK(clk), .Q(
        regs[254]) );
  EDQV2_8TH40 regs_reg_24__29_ ( .D(wdata[29]), .E(n1247), .CK(clk), .Q(
        regs[253]) );
  EDQV2_8TH40 regs_reg_24__28_ ( .D(wdata[28]), .E(n1247), .CK(clk), .Q(
        regs[252]) );
  EDQV2_8TH40 regs_reg_24__27_ ( .D(wdata[27]), .E(n1247), .CK(clk), .Q(
        regs[251]) );
  EDQV2_8TH40 regs_reg_24__26_ ( .D(wdata[26]), .E(n1247), .CK(clk), .Q(
        regs[250]) );
  EDQV2_8TH40 regs_reg_24__25_ ( .D(wdata[25]), .E(n1247), .CK(clk), .Q(
        regs[249]) );
  EDQV2_8TH40 regs_reg_24__24_ ( .D(wdata[24]), .E(n1247), .CK(clk), .Q(
        regs[248]) );
  EDQV2_8TH40 regs_reg_24__23_ ( .D(wdata[23]), .E(n1247), .CK(clk), .Q(
        regs[247]) );
  EDQV2_8TH40 regs_reg_24__22_ ( .D(wdata[22]), .E(n1247), .CK(clk), .Q(
        regs[246]) );
  EDQV2_8TH40 regs_reg_24__21_ ( .D(wdata[21]), .E(n1247), .CK(clk), .Q(
        regs[245]) );
  EDQV2_8TH40 regs_reg_24__20_ ( .D(wdata[20]), .E(n1247), .CK(clk), .Q(
        regs[244]) );
  EDQV2_8TH40 regs_reg_24__19_ ( .D(wdata[19]), .E(n1247), .CK(clk), .Q(
        regs[243]) );
  EDQV2_8TH40 regs_reg_24__18_ ( .D(wdata[18]), .E(n1247), .CK(clk), .Q(
        regs[242]) );
  EDQV2_8TH40 regs_reg_24__17_ ( .D(wdata[17]), .E(n1247), .CK(clk), .Q(
        regs[241]) );
  EDQV2_8TH40 regs_reg_24__16_ ( .D(wdata[16]), .E(n1247), .CK(clk), .Q(
        regs[240]) );
  EDQV2_8TH40 regs_reg_24__15_ ( .D(wdata[15]), .E(n1247), .CK(clk), .Q(
        regs[239]) );
  EDQV2_8TH40 regs_reg_24__14_ ( .D(wdata[14]), .E(n1247), .CK(clk), .Q(
        regs[238]) );
  EDQV2_8TH40 regs_reg_24__13_ ( .D(wdata[13]), .E(n1247), .CK(clk), .Q(
        regs[237]) );
  EDQV2_8TH40 regs_reg_24__12_ ( .D(wdata[12]), .E(n1247), .CK(clk), .Q(
        regs[236]) );
  EDQV2_8TH40 regs_reg_24__11_ ( .D(wdata[11]), .E(n1247), .CK(clk), .Q(
        regs[235]) );
  EDQV2_8TH40 regs_reg_24__10_ ( .D(wdata[10]), .E(n1247), .CK(clk), .Q(
        regs[234]) );
  EDQV2_8TH40 regs_reg_24__9_ ( .D(wdata[9]), .E(n1247), .CK(clk), .Q(
        regs[233]) );
  EDQV2_8TH40 regs_reg_24__8_ ( .D(wdata[8]), .E(n1247), .CK(clk), .Q(
        regs[232]) );
  EDQV2_8TH40 regs_reg_24__7_ ( .D(wdata[7]), .E(n1247), .CK(clk), .Q(
        regs[231]) );
  EDQV2_8TH40 regs_reg_24__6_ ( .D(wdata[6]), .E(n1247), .CK(clk), .Q(
        regs[230]) );
  EDQV2_8TH40 regs_reg_24__5_ ( .D(wdata[5]), .E(n1247), .CK(clk), .Q(
        regs[229]) );
  EDQV2_8TH40 regs_reg_24__4_ ( .D(wdata[4]), .E(n1247), .CK(clk), .Q(
        regs[228]) );
  EDQV2_8TH40 regs_reg_24__3_ ( .D(wdata[3]), .E(n1247), .CK(clk), .Q(
        regs[227]) );
  EDQV2_8TH40 regs_reg_24__2_ ( .D(wdata[2]), .E(n1247), .CK(clk), .Q(
        regs[226]) );
  EDQV2_8TH40 regs_reg_24__1_ ( .D(wdata[1]), .E(n1247), .CK(clk), .Q(
        regs[225]) );
  EDQV2_8TH40 regs_reg_24__0_ ( .D(wdata[0]), .E(n1247), .CK(clk), .Q(
        regs[224]) );
  EDQV2_8TH40 regs_reg_28__31_ ( .D(wdata[31]), .E(n1250), .CK(clk), .Q(
        regs[127]) );
  EDQV2_8TH40 regs_reg_28__30_ ( .D(wdata[30]), .E(n1250), .CK(clk), .Q(
        regs[126]) );
  EDQV2_8TH40 regs_reg_28__29_ ( .D(wdata[29]), .E(n1250), .CK(clk), .Q(
        regs[125]) );
  EDQV2_8TH40 regs_reg_28__28_ ( .D(wdata[28]), .E(n1250), .CK(clk), .Q(
        regs[124]) );
  EDQV2_8TH40 regs_reg_28__27_ ( .D(wdata[27]), .E(n1250), .CK(clk), .Q(
        regs[123]) );
  EDQV2_8TH40 regs_reg_28__26_ ( .D(wdata[26]), .E(n1250), .CK(clk), .Q(
        regs[122]) );
  EDQV2_8TH40 regs_reg_28__25_ ( .D(wdata[25]), .E(n1250), .CK(clk), .Q(
        regs[121]) );
  EDQV2_8TH40 regs_reg_28__24_ ( .D(wdata[24]), .E(n1250), .CK(clk), .Q(
        regs[120]) );
  EDQV2_8TH40 regs_reg_28__23_ ( .D(wdata[23]), .E(n1250), .CK(clk), .Q(
        regs[119]) );
  EDQV2_8TH40 regs_reg_28__22_ ( .D(wdata[22]), .E(n1250), .CK(clk), .Q(
        regs[118]) );
  EDQV2_8TH40 regs_reg_28__21_ ( .D(wdata[21]), .E(n1250), .CK(clk), .Q(
        regs[117]) );
  EDQV2_8TH40 regs_reg_28__20_ ( .D(wdata[20]), .E(n1250), .CK(clk), .Q(
        regs[116]) );
  EDQV2_8TH40 regs_reg_28__19_ ( .D(wdata[19]), .E(n1250), .CK(clk), .Q(
        regs[115]) );
  EDQV2_8TH40 regs_reg_28__18_ ( .D(wdata[18]), .E(n1250), .CK(clk), .Q(
        regs[114]) );
  EDQV2_8TH40 regs_reg_28__17_ ( .D(wdata[17]), .E(n1250), .CK(clk), .Q(
        regs[113]) );
  EDQV2_8TH40 regs_reg_28__16_ ( .D(wdata[16]), .E(n1250), .CK(clk), .Q(
        regs[112]) );
  EDQV2_8TH40 regs_reg_28__15_ ( .D(wdata[15]), .E(n1250), .CK(clk), .Q(
        regs[111]) );
  EDQV2_8TH40 regs_reg_28__14_ ( .D(wdata[14]), .E(n1250), .CK(clk), .Q(
        regs[110]) );
  EDQV2_8TH40 regs_reg_28__13_ ( .D(wdata[13]), .E(n1250), .CK(clk), .Q(
        regs[109]) );
  EDQV2_8TH40 regs_reg_28__12_ ( .D(wdata[12]), .E(n1250), .CK(clk), .Q(
        regs[108]) );
  EDQV2_8TH40 regs_reg_28__11_ ( .D(wdata[11]), .E(n1250), .CK(clk), .Q(
        regs[107]) );
  EDQV2_8TH40 regs_reg_28__10_ ( .D(wdata[10]), .E(n1250), .CK(clk), .Q(
        regs[106]) );
  EDQV2_8TH40 regs_reg_28__9_ ( .D(wdata[9]), .E(n1250), .CK(clk), .Q(
        regs[105]) );
  EDQV2_8TH40 regs_reg_28__8_ ( .D(wdata[8]), .E(n1250), .CK(clk), .Q(
        regs[104]) );
  EDQV2_8TH40 regs_reg_28__7_ ( .D(wdata[7]), .E(n1250), .CK(clk), .Q(
        regs[103]) );
  EDQV2_8TH40 regs_reg_28__6_ ( .D(wdata[6]), .E(n1250), .CK(clk), .Q(
        regs[102]) );
  EDQV2_8TH40 regs_reg_28__5_ ( .D(wdata[5]), .E(n1250), .CK(clk), .Q(
        regs[101]) );
  EDQV2_8TH40 regs_reg_28__4_ ( .D(wdata[4]), .E(n1250), .CK(clk), .Q(
        regs[100]) );
  EDQV2_8TH40 regs_reg_28__3_ ( .D(wdata[3]), .E(n1250), .CK(clk), .Q(regs[99]) );
  EDQV2_8TH40 regs_reg_28__2_ ( .D(wdata[2]), .E(n1250), .CK(clk), .Q(regs[98]) );
  EDQV2_8TH40 regs_reg_28__1_ ( .D(wdata[1]), .E(n1250), .CK(clk), .Q(regs[97]) );
  EDQV2_8TH40 regs_reg_28__0_ ( .D(wdata[0]), .E(n1250), .CK(clk), .Q(regs[96]) );
  EDQV2_8TH40 regs_reg_1__31_ ( .D(wdata[31]), .E(n1233), .CK(clk), .Q(
        regs[991]) );
  EDQV2_8TH40 regs_reg_1__30_ ( .D(wdata[30]), .E(n1233), .CK(clk), .Q(
        regs[990]) );
  EDQV2_8TH40 regs_reg_1__29_ ( .D(wdata[29]), .E(n1233), .CK(clk), .Q(
        regs[989]) );
  EDQV2_8TH40 regs_reg_1__28_ ( .D(wdata[28]), .E(n1233), .CK(clk), .Q(
        regs[988]) );
  EDQV2_8TH40 regs_reg_1__27_ ( .D(wdata[27]), .E(n1233), .CK(clk), .Q(
        regs[987]) );
  EDQV2_8TH40 regs_reg_1__26_ ( .D(wdata[26]), .E(n1233), .CK(clk), .Q(
        regs[986]) );
  EDQV2_8TH40 regs_reg_1__25_ ( .D(wdata[25]), .E(n1233), .CK(clk), .Q(
        regs[985]) );
  EDQV2_8TH40 regs_reg_1__24_ ( .D(wdata[24]), .E(n1233), .CK(clk), .Q(
        regs[984]) );
  EDQV2_8TH40 regs_reg_1__23_ ( .D(wdata[23]), .E(n1233), .CK(clk), .Q(
        regs[983]) );
  EDQV2_8TH40 regs_reg_1__22_ ( .D(wdata[22]), .E(n1233), .CK(clk), .Q(
        regs[982]) );
  EDQV2_8TH40 regs_reg_1__21_ ( .D(wdata[21]), .E(n1233), .CK(clk), .Q(
        regs[981]) );
  EDQV2_8TH40 regs_reg_1__20_ ( .D(wdata[20]), .E(n1233), .CK(clk), .Q(
        regs[980]) );
  EDQV2_8TH40 regs_reg_1__19_ ( .D(wdata[19]), .E(n1233), .CK(clk), .Q(
        regs[979]) );
  EDQV2_8TH40 regs_reg_1__18_ ( .D(wdata[18]), .E(n1233), .CK(clk), .Q(
        regs[978]) );
  EDQV2_8TH40 regs_reg_1__17_ ( .D(wdata[17]), .E(n1233), .CK(clk), .Q(
        regs[977]) );
  EDQV2_8TH40 regs_reg_1__16_ ( .D(wdata[16]), .E(n1233), .CK(clk), .Q(
        regs[976]) );
  EDQV2_8TH40 regs_reg_1__15_ ( .D(wdata[15]), .E(n1233), .CK(clk), .Q(
        regs[975]) );
  EDQV2_8TH40 regs_reg_1__14_ ( .D(wdata[14]), .E(n1233), .CK(clk), .Q(
        regs[974]) );
  EDQV2_8TH40 regs_reg_1__13_ ( .D(wdata[13]), .E(n1233), .CK(clk), .Q(
        regs[973]) );
  EDQV2_8TH40 regs_reg_1__12_ ( .D(wdata[12]), .E(n1233), .CK(clk), .Q(
        regs[972]) );
  EDQV2_8TH40 regs_reg_1__11_ ( .D(wdata[11]), .E(n1233), .CK(clk), .Q(
        regs[971]) );
  EDQV2_8TH40 regs_reg_1__10_ ( .D(wdata[10]), .E(n1233), .CK(clk), .Q(
        regs[970]) );
  EDQV2_8TH40 regs_reg_1__9_ ( .D(wdata[9]), .E(n1233), .CK(clk), .Q(regs[969]) );
  EDQV2_8TH40 regs_reg_1__8_ ( .D(wdata[8]), .E(n1233), .CK(clk), .Q(regs[968]) );
  EDQV2_8TH40 regs_reg_1__7_ ( .D(wdata[7]), .E(n1233), .CK(clk), .Q(regs[967]) );
  EDQV2_8TH40 regs_reg_1__6_ ( .D(wdata[6]), .E(n1233), .CK(clk), .Q(regs[966]) );
  EDQV2_8TH40 regs_reg_1__5_ ( .D(wdata[5]), .E(n1233), .CK(clk), .Q(regs[965]) );
  EDQV2_8TH40 regs_reg_1__4_ ( .D(wdata[4]), .E(n1233), .CK(clk), .Q(regs[964]) );
  EDQV2_8TH40 regs_reg_1__3_ ( .D(wdata[3]), .E(n1233), .CK(clk), .Q(regs[963]) );
  EDQV2_8TH40 regs_reg_1__2_ ( .D(wdata[2]), .E(n1233), .CK(clk), .Q(regs[962]) );
  EDQV2_8TH40 regs_reg_1__1_ ( .D(wdata[1]), .E(n1233), .CK(clk), .Q(regs[961]) );
  EDQV2_8TH40 regs_reg_1__0_ ( .D(wdata[0]), .E(n1233), .CK(clk), .Q(regs[960]) );
  EDQV2_8TH40 regs_reg_9__31_ ( .D(wdata[31]), .E(n1237), .CK(clk), .Q(
        regs[735]) );
  EDQV2_8TH40 regs_reg_9__30_ ( .D(wdata[30]), .E(n1237), .CK(clk), .Q(
        regs[734]) );
  EDQV2_8TH40 regs_reg_9__29_ ( .D(wdata[29]), .E(n1237), .CK(clk), .Q(
        regs[733]) );
  EDQV2_8TH40 regs_reg_9__28_ ( .D(wdata[28]), .E(n1237), .CK(clk), .Q(
        regs[732]) );
  EDQV2_8TH40 regs_reg_9__27_ ( .D(wdata[27]), .E(n1237), .CK(clk), .Q(
        regs[731]) );
  EDQV2_8TH40 regs_reg_9__26_ ( .D(wdata[26]), .E(n1237), .CK(clk), .Q(
        regs[730]) );
  EDQV2_8TH40 regs_reg_9__25_ ( .D(wdata[25]), .E(n1237), .CK(clk), .Q(
        regs[729]) );
  EDQV2_8TH40 regs_reg_9__24_ ( .D(wdata[24]), .E(n1237), .CK(clk), .Q(
        regs[728]) );
  EDQV2_8TH40 regs_reg_9__23_ ( .D(wdata[23]), .E(n1237), .CK(clk), .Q(
        regs[727]) );
  EDQV2_8TH40 regs_reg_9__22_ ( .D(wdata[22]), .E(n1237), .CK(clk), .Q(
        regs[726]) );
  EDQV2_8TH40 regs_reg_9__21_ ( .D(wdata[21]), .E(n1237), .CK(clk), .Q(
        regs[725]) );
  EDQV2_8TH40 regs_reg_9__20_ ( .D(wdata[20]), .E(n1237), .CK(clk), .Q(
        regs[724]) );
  EDQV2_8TH40 regs_reg_9__19_ ( .D(wdata[19]), .E(n1237), .CK(clk), .Q(
        regs[723]) );
  EDQV2_8TH40 regs_reg_9__18_ ( .D(wdata[18]), .E(n1237), .CK(clk), .Q(
        regs[722]) );
  EDQV2_8TH40 regs_reg_9__17_ ( .D(wdata[17]), .E(n1237), .CK(clk), .Q(
        regs[721]) );
  EDQV2_8TH40 regs_reg_9__16_ ( .D(wdata[16]), .E(n1237), .CK(clk), .Q(
        regs[720]) );
  EDQV2_8TH40 regs_reg_9__15_ ( .D(wdata[15]), .E(n1237), .CK(clk), .Q(
        regs[719]) );
  EDQV2_8TH40 regs_reg_9__14_ ( .D(wdata[14]), .E(n1237), .CK(clk), .Q(
        regs[718]) );
  EDQV2_8TH40 regs_reg_9__13_ ( .D(wdata[13]), .E(n1237), .CK(clk), .Q(
        regs[717]) );
  EDQV2_8TH40 regs_reg_9__12_ ( .D(wdata[12]), .E(n1237), .CK(clk), .Q(
        regs[716]) );
  EDQV2_8TH40 regs_reg_9__11_ ( .D(wdata[11]), .E(n1237), .CK(clk), .Q(
        regs[715]) );
  EDQV2_8TH40 regs_reg_9__10_ ( .D(wdata[10]), .E(n1237), .CK(clk), .Q(
        regs[714]) );
  EDQV2_8TH40 regs_reg_9__9_ ( .D(wdata[9]), .E(n1237), .CK(clk), .Q(regs[713]) );
  EDQV2_8TH40 regs_reg_9__8_ ( .D(wdata[8]), .E(n1237), .CK(clk), .Q(regs[712]) );
  EDQV2_8TH40 regs_reg_9__7_ ( .D(wdata[7]), .E(n1237), .CK(clk), .Q(regs[711]) );
  EDQV2_8TH40 regs_reg_9__6_ ( .D(wdata[6]), .E(n1237), .CK(clk), .Q(regs[710]) );
  EDQV2_8TH40 regs_reg_9__5_ ( .D(wdata[5]), .E(n1237), .CK(clk), .Q(regs[709]) );
  EDQV2_8TH40 regs_reg_9__4_ ( .D(wdata[4]), .E(n1237), .CK(clk), .Q(regs[708]) );
  EDQV2_8TH40 regs_reg_9__3_ ( .D(wdata[3]), .E(n1237), .CK(clk), .Q(regs[707]) );
  EDQV2_8TH40 regs_reg_9__2_ ( .D(wdata[2]), .E(n1237), .CK(clk), .Q(regs[706]) );
  EDQV2_8TH40 regs_reg_9__1_ ( .D(wdata[1]), .E(n1237), .CK(clk), .Q(regs[705]) );
  EDQV2_8TH40 regs_reg_9__0_ ( .D(wdata[0]), .E(n1237), .CK(clk), .Q(regs[704]) );
  EDQV2_8TH40 regs_reg_17__31_ ( .D(wdata[31]), .E(n1241), .CK(clk), .Q(
        regs[479]) );
  EDQV2_8TH40 regs_reg_17__30_ ( .D(wdata[30]), .E(n1241), .CK(clk), .Q(
        regs[478]) );
  EDQV2_8TH40 regs_reg_17__29_ ( .D(wdata[29]), .E(n1241), .CK(clk), .Q(
        regs[477]) );
  EDQV2_8TH40 regs_reg_17__28_ ( .D(wdata[28]), .E(n1241), .CK(clk), .Q(
        regs[476]) );
  EDQV2_8TH40 regs_reg_17__27_ ( .D(wdata[27]), .E(n1241), .CK(clk), .Q(
        regs[475]) );
  EDQV2_8TH40 regs_reg_17__26_ ( .D(wdata[26]), .E(n1241), .CK(clk), .Q(
        regs[474]) );
  EDQV2_8TH40 regs_reg_17__25_ ( .D(wdata[25]), .E(n1241), .CK(clk), .Q(
        regs[473]) );
  EDQV2_8TH40 regs_reg_17__24_ ( .D(wdata[24]), .E(n1241), .CK(clk), .Q(
        regs[472]) );
  EDQV2_8TH40 regs_reg_17__23_ ( .D(wdata[23]), .E(n1241), .CK(clk), .Q(
        regs[471]) );
  EDQV2_8TH40 regs_reg_17__22_ ( .D(wdata[22]), .E(n1241), .CK(clk), .Q(
        regs[470]) );
  EDQV2_8TH40 regs_reg_17__21_ ( .D(wdata[21]), .E(n1241), .CK(clk), .Q(
        regs[469]) );
  EDQV2_8TH40 regs_reg_17__20_ ( .D(wdata[20]), .E(n1241), .CK(clk), .Q(
        regs[468]) );
  EDQV2_8TH40 regs_reg_17__19_ ( .D(wdata[19]), .E(n1241), .CK(clk), .Q(
        regs[467]) );
  EDQV2_8TH40 regs_reg_17__18_ ( .D(wdata[18]), .E(n1241), .CK(clk), .Q(
        regs[466]) );
  EDQV2_8TH40 regs_reg_17__17_ ( .D(wdata[17]), .E(n1241), .CK(clk), .Q(
        regs[465]) );
  EDQV2_8TH40 regs_reg_17__16_ ( .D(wdata[16]), .E(n1241), .CK(clk), .Q(
        regs[464]) );
  EDQV2_8TH40 regs_reg_17__15_ ( .D(wdata[15]), .E(n1241), .CK(clk), .Q(
        regs[463]) );
  EDQV2_8TH40 regs_reg_17__14_ ( .D(wdata[14]), .E(n1241), .CK(clk), .Q(
        regs[462]) );
  EDQV2_8TH40 regs_reg_17__13_ ( .D(wdata[13]), .E(n1241), .CK(clk), .Q(
        regs[461]) );
  EDQV2_8TH40 regs_reg_17__12_ ( .D(wdata[12]), .E(n1241), .CK(clk), .Q(
        regs[460]) );
  EDQV2_8TH40 regs_reg_17__11_ ( .D(wdata[11]), .E(n1241), .CK(clk), .Q(
        regs[459]) );
  EDQV2_8TH40 regs_reg_17__10_ ( .D(wdata[10]), .E(n1241), .CK(clk), .Q(
        regs[458]) );
  EDQV2_8TH40 regs_reg_17__9_ ( .D(wdata[9]), .E(n1241), .CK(clk), .Q(
        regs[457]) );
  EDQV2_8TH40 regs_reg_17__8_ ( .D(wdata[8]), .E(n1241), .CK(clk), .Q(
        regs[456]) );
  EDQV2_8TH40 regs_reg_17__7_ ( .D(wdata[7]), .E(n1241), .CK(clk), .Q(
        regs[455]) );
  EDQV2_8TH40 regs_reg_17__6_ ( .D(wdata[6]), .E(n1241), .CK(clk), .Q(
        regs[454]) );
  EDQV2_8TH40 regs_reg_17__5_ ( .D(wdata[5]), .E(n1241), .CK(clk), .Q(
        regs[453]) );
  EDQV2_8TH40 regs_reg_17__4_ ( .D(wdata[4]), .E(n1241), .CK(clk), .Q(
        regs[452]) );
  EDQV2_8TH40 regs_reg_17__3_ ( .D(wdata[3]), .E(n1241), .CK(clk), .Q(
        regs[451]) );
  EDQV2_8TH40 regs_reg_17__2_ ( .D(wdata[2]), .E(n1241), .CK(clk), .Q(
        regs[450]) );
  EDQV2_8TH40 regs_reg_17__1_ ( .D(wdata[1]), .E(n1241), .CK(clk), .Q(
        regs[449]) );
  EDQV2_8TH40 regs_reg_17__0_ ( .D(wdata[0]), .E(n1241), .CK(clk), .Q(
        regs[448]) );
  EDQV2_8TH40 regs_reg_21__31_ ( .D(wdata[31]), .E(n1245), .CK(clk), .Q(
        regs[351]) );
  EDQV2_8TH40 regs_reg_21__30_ ( .D(wdata[30]), .E(n1245), .CK(clk), .Q(
        regs[350]) );
  EDQV2_8TH40 regs_reg_21__29_ ( .D(wdata[29]), .E(n1245), .CK(clk), .Q(
        regs[349]) );
  EDQV2_8TH40 regs_reg_21__28_ ( .D(wdata[28]), .E(n1245), .CK(clk), .Q(
        regs[348]) );
  EDQV2_8TH40 regs_reg_21__27_ ( .D(wdata[27]), .E(n1245), .CK(clk), .Q(
        regs[347]) );
  EDQV2_8TH40 regs_reg_21__26_ ( .D(wdata[26]), .E(n1245), .CK(clk), .Q(
        regs[346]) );
  EDQV2_8TH40 regs_reg_21__25_ ( .D(wdata[25]), .E(n1245), .CK(clk), .Q(
        regs[345]) );
  EDQV2_8TH40 regs_reg_21__24_ ( .D(wdata[24]), .E(n1245), .CK(clk), .Q(
        regs[344]) );
  EDQV2_8TH40 regs_reg_21__23_ ( .D(wdata[23]), .E(n1245), .CK(clk), .Q(
        regs[343]) );
  EDQV2_8TH40 regs_reg_21__22_ ( .D(wdata[22]), .E(n1245), .CK(clk), .Q(
        regs[342]) );
  EDQV2_8TH40 regs_reg_21__21_ ( .D(wdata[21]), .E(n1245), .CK(clk), .Q(
        regs[341]) );
  EDQV2_8TH40 regs_reg_21__20_ ( .D(wdata[20]), .E(n1245), .CK(clk), .Q(
        regs[340]) );
  EDQV2_8TH40 regs_reg_21__19_ ( .D(wdata[19]), .E(n1245), .CK(clk), .Q(
        regs[339]) );
  EDQV2_8TH40 regs_reg_21__18_ ( .D(wdata[18]), .E(n1245), .CK(clk), .Q(
        regs[338]) );
  EDQV2_8TH40 regs_reg_21__17_ ( .D(wdata[17]), .E(n1245), .CK(clk), .Q(
        regs[337]) );
  EDQV2_8TH40 regs_reg_21__16_ ( .D(wdata[16]), .E(n1245), .CK(clk), .Q(
        regs[336]) );
  EDQV2_8TH40 regs_reg_21__15_ ( .D(wdata[15]), .E(n1245), .CK(clk), .Q(
        regs[335]) );
  EDQV2_8TH40 regs_reg_21__14_ ( .D(wdata[14]), .E(n1245), .CK(clk), .Q(
        regs[334]) );
  EDQV2_8TH40 regs_reg_21__13_ ( .D(wdata[13]), .E(n1245), .CK(clk), .Q(
        regs[333]) );
  EDQV2_8TH40 regs_reg_21__12_ ( .D(wdata[12]), .E(n1245), .CK(clk), .Q(
        regs[332]) );
  EDQV2_8TH40 regs_reg_21__11_ ( .D(wdata[11]), .E(n1245), .CK(clk), .Q(
        regs[331]) );
  EDQV2_8TH40 regs_reg_21__10_ ( .D(wdata[10]), .E(n1245), .CK(clk), .Q(
        regs[330]) );
  EDQV2_8TH40 regs_reg_21__9_ ( .D(wdata[9]), .E(n1245), .CK(clk), .Q(
        regs[329]) );
  EDQV2_8TH40 regs_reg_21__8_ ( .D(wdata[8]), .E(n1245), .CK(clk), .Q(
        regs[328]) );
  EDQV2_8TH40 regs_reg_21__7_ ( .D(wdata[7]), .E(n1245), .CK(clk), .Q(
        regs[327]) );
  EDQV2_8TH40 regs_reg_21__6_ ( .D(wdata[6]), .E(n1245), .CK(clk), .Q(
        regs[326]) );
  EDQV2_8TH40 regs_reg_21__5_ ( .D(wdata[5]), .E(n1245), .CK(clk), .Q(
        regs[325]) );
  EDQV2_8TH40 regs_reg_21__4_ ( .D(wdata[4]), .E(n1245), .CK(clk), .Q(
        regs[324]) );
  EDQV2_8TH40 regs_reg_21__3_ ( .D(wdata[3]), .E(n1245), .CK(clk), .Q(
        regs[323]) );
  EDQV2_8TH40 regs_reg_21__2_ ( .D(wdata[2]), .E(n1245), .CK(clk), .Q(
        regs[322]) );
  EDQV2_8TH40 regs_reg_21__1_ ( .D(wdata[1]), .E(n1245), .CK(clk), .Q(
        regs[321]) );
  EDQV2_8TH40 regs_reg_21__0_ ( .D(wdata[0]), .E(n1245), .CK(clk), .Q(
        regs[320]) );
  EDQV2_8TH40 regs_reg_25__31_ ( .D(wdata[31]), .E(n1248), .CK(clk), .Q(
        regs[223]) );
  EDQV2_8TH40 regs_reg_25__30_ ( .D(wdata[30]), .E(n1248), .CK(clk), .Q(
        regs[222]) );
  EDQV2_8TH40 regs_reg_25__29_ ( .D(wdata[29]), .E(n1248), .CK(clk), .Q(
        regs[221]) );
  EDQV2_8TH40 regs_reg_25__28_ ( .D(wdata[28]), .E(n1248), .CK(clk), .Q(
        regs[220]) );
  EDQV2_8TH40 regs_reg_25__27_ ( .D(wdata[27]), .E(n1248), .CK(clk), .Q(
        regs[219]) );
  EDQV2_8TH40 regs_reg_25__26_ ( .D(wdata[26]), .E(n1248), .CK(clk), .Q(
        regs[218]) );
  EDQV2_8TH40 regs_reg_25__25_ ( .D(wdata[25]), .E(n1248), .CK(clk), .Q(
        regs[217]) );
  EDQV2_8TH40 regs_reg_25__24_ ( .D(wdata[24]), .E(n1248), .CK(clk), .Q(
        regs[216]) );
  EDQV2_8TH40 regs_reg_25__23_ ( .D(wdata[23]), .E(n1248), .CK(clk), .Q(
        regs[215]) );
  EDQV2_8TH40 regs_reg_25__22_ ( .D(wdata[22]), .E(n1248), .CK(clk), .Q(
        regs[214]) );
  EDQV2_8TH40 regs_reg_25__21_ ( .D(wdata[21]), .E(n1248), .CK(clk), .Q(
        regs[213]) );
  EDQV2_8TH40 regs_reg_25__20_ ( .D(wdata[20]), .E(n1248), .CK(clk), .Q(
        regs[212]) );
  EDQV2_8TH40 regs_reg_25__19_ ( .D(wdata[19]), .E(n1248), .CK(clk), .Q(
        regs[211]) );
  EDQV2_8TH40 regs_reg_25__18_ ( .D(wdata[18]), .E(n1248), .CK(clk), .Q(
        regs[210]) );
  EDQV2_8TH40 regs_reg_25__17_ ( .D(wdata[17]), .E(n1248), .CK(clk), .Q(
        regs[209]) );
  EDQV2_8TH40 regs_reg_25__16_ ( .D(wdata[16]), .E(n1248), .CK(clk), .Q(
        regs[208]) );
  EDQV2_8TH40 regs_reg_25__15_ ( .D(wdata[15]), .E(n1248), .CK(clk), .Q(
        regs[207]) );
  EDQV2_8TH40 regs_reg_25__14_ ( .D(wdata[14]), .E(n1248), .CK(clk), .Q(
        regs[206]) );
  EDQV2_8TH40 regs_reg_25__13_ ( .D(wdata[13]), .E(n1248), .CK(clk), .Q(
        regs[205]) );
  EDQV2_8TH40 regs_reg_25__12_ ( .D(wdata[12]), .E(n1248), .CK(clk), .Q(
        regs[204]) );
  EDQV2_8TH40 regs_reg_25__11_ ( .D(wdata[11]), .E(n1248), .CK(clk), .Q(
        regs[203]) );
  EDQV2_8TH40 regs_reg_25__10_ ( .D(wdata[10]), .E(n1248), .CK(clk), .Q(
        regs[202]) );
  EDQV2_8TH40 regs_reg_25__9_ ( .D(wdata[9]), .E(n1248), .CK(clk), .Q(
        regs[201]) );
  EDQV2_8TH40 regs_reg_25__8_ ( .D(wdata[8]), .E(n1248), .CK(clk), .Q(
        regs[200]) );
  EDQV2_8TH40 regs_reg_25__7_ ( .D(wdata[7]), .E(n1248), .CK(clk), .Q(
        regs[199]) );
  EDQV2_8TH40 regs_reg_25__6_ ( .D(wdata[6]), .E(n1248), .CK(clk), .Q(
        regs[198]) );
  EDQV2_8TH40 regs_reg_25__5_ ( .D(wdata[5]), .E(n1248), .CK(clk), .Q(
        regs[197]) );
  EDQV2_8TH40 regs_reg_25__4_ ( .D(wdata[4]), .E(n1248), .CK(clk), .Q(
        regs[196]) );
  EDQV2_8TH40 regs_reg_25__3_ ( .D(wdata[3]), .E(n1248), .CK(clk), .Q(
        regs[195]) );
  EDQV2_8TH40 regs_reg_25__2_ ( .D(wdata[2]), .E(n1248), .CK(clk), .Q(
        regs[194]) );
  EDQV2_8TH40 regs_reg_25__1_ ( .D(wdata[1]), .E(n1248), .CK(clk), .Q(
        regs[193]) );
  EDQV2_8TH40 regs_reg_25__0_ ( .D(wdata[0]), .E(n1248), .CK(clk), .Q(
        regs[192]) );
  DQV2_8TH40 regs_reg_0__31_ ( .D(regs[1023]), .CK(clk), .Q(regs[1023]) );
  DQV2_8TH40 regs_reg_0__30_ ( .D(regs[1022]), .CK(clk), .Q(regs[1022]) );
  DQV2_8TH40 regs_reg_0__29_ ( .D(regs[1021]), .CK(clk), .Q(regs[1021]) );
  DQV2_8TH40 regs_reg_0__28_ ( .D(regs[1020]), .CK(clk), .Q(regs[1020]) );
  DQV2_8TH40 regs_reg_0__27_ ( .D(regs[1019]), .CK(clk), .Q(regs[1019]) );
  DQV2_8TH40 regs_reg_0__26_ ( .D(regs[1018]), .CK(clk), .Q(regs[1018]) );
  DQV2_8TH40 regs_reg_0__25_ ( .D(regs[1017]), .CK(clk), .Q(regs[1017]) );
  DQV2_8TH40 regs_reg_0__24_ ( .D(regs[1016]), .CK(clk), .Q(regs[1016]) );
  DQV2_8TH40 regs_reg_0__23_ ( .D(regs[1015]), .CK(clk), .Q(regs[1015]) );
  DQV2_8TH40 regs_reg_0__22_ ( .D(regs[1014]), .CK(clk), .Q(regs[1014]) );
  DQV2_8TH40 regs_reg_0__21_ ( .D(regs[1013]), .CK(clk), .Q(regs[1013]) );
  DQV2_8TH40 regs_reg_0__20_ ( .D(regs[1012]), .CK(clk), .Q(regs[1012]) );
  DQV2_8TH40 regs_reg_0__19_ ( .D(regs[1011]), .CK(clk), .Q(regs[1011]) );
  DQV2_8TH40 regs_reg_0__18_ ( .D(regs[1010]), .CK(clk), .Q(regs[1010]) );
  DQV2_8TH40 regs_reg_0__17_ ( .D(regs[1009]), .CK(clk), .Q(regs[1009]) );
  DQV2_8TH40 regs_reg_0__16_ ( .D(regs[1008]), .CK(clk), .Q(regs[1008]) );
  DQV2_8TH40 regs_reg_0__15_ ( .D(regs[1007]), .CK(clk), .Q(regs[1007]) );
  DQV2_8TH40 regs_reg_0__14_ ( .D(regs[1006]), .CK(clk), .Q(regs[1006]) );
  DQV2_8TH40 regs_reg_0__13_ ( .D(regs[1005]), .CK(clk), .Q(regs[1005]) );
  DQV2_8TH40 regs_reg_0__12_ ( .D(regs[1004]), .CK(clk), .Q(regs[1004]) );
  DQV2_8TH40 regs_reg_0__11_ ( .D(regs[1003]), .CK(clk), .Q(regs[1003]) );
  DQV2_8TH40 regs_reg_0__10_ ( .D(regs[1002]), .CK(clk), .Q(regs[1002]) );
  DQV2_8TH40 regs_reg_0__9_ ( .D(regs[1001]), .CK(clk), .Q(regs[1001]) );
  DQV2_8TH40 regs_reg_0__8_ ( .D(regs[1000]), .CK(clk), .Q(regs[1000]) );
  DQV2_8TH40 regs_reg_0__7_ ( .D(regs[999]), .CK(clk), .Q(regs[999]) );
  DQV2_8TH40 regs_reg_0__6_ ( .D(regs[998]), .CK(clk), .Q(regs[998]) );
  DQV2_8TH40 regs_reg_0__5_ ( .D(regs[997]), .CK(clk), .Q(regs[997]) );
  DQV2_8TH40 regs_reg_0__4_ ( .D(regs[996]), .CK(clk), .Q(regs[996]) );
  DQV2_8TH40 regs_reg_0__3_ ( .D(regs[995]), .CK(clk), .Q(regs[995]) );
  DQV2_8TH40 regs_reg_0__2_ ( .D(regs[994]), .CK(clk), .Q(regs[994]) );
  DQV2_8TH40 regs_reg_0__1_ ( .D(regs[993]), .CK(clk), .Q(regs[993]) );
  DQV2_8TH40 regs_reg_0__0_ ( .D(regs[992]), .CK(clk), .Q(regs[992]) );
  I2NOR4V2_8TH40 U2 ( .A1(re1), .A2(n1195), .B1(n1196), .B2(rst), .ZN(n1194)
         );
  IOA22V4_8TH40 U3 ( .B1(n1154), .B2(n1193), .A1(N121), .A2(n1194), .ZN(
        rdata1[5]) );
  CKMUX2V8_8TH40 U4 ( .I0(n567), .I1(n562), .S(raddr1[4]), .Z(N121) );
  CKMUX2V8_8TH40 U5 ( .I0(n577), .I1(n572), .S(raddr1[4]), .Z(N120) );
  CKMUX2V8_8TH40 U6 ( .I0(n587), .I1(n582), .S(raddr1[4]), .Z(N119) );
  CKMUX2V8_8TH40 U7 ( .I0(n597), .I1(n592), .S(raddr1[4]), .Z(N118) );
  CKMUX2V8_8TH40 U8 ( .I0(n607), .I1(n602), .S(raddr1[4]), .Z(N117) );
  CKMUX2V8_8TH40 U9 ( .I0(n617), .I1(n612), .S(raddr1[4]), .Z(N116) );
  CKMUX2V8_8TH40 U10 ( .I0(n627), .I1(n622), .S(raddr1[4]), .Z(N115) );
  CKMUX2V8_8TH40 U11 ( .I0(n637), .I1(n632), .S(raddr1[4]), .Z(N114) );
  CKMUX2V8_8TH40 U12 ( .I0(n647), .I1(n642), .S(raddr1[4]), .Z(N113) );
  CKMUX2V8_8TH40 U13 ( .I0(n657), .I1(n652), .S(raddr1[4]), .Z(N112) );
  CKMUX2V8_8TH40 U14 ( .I0(n667), .I1(n662), .S(raddr1[4]), .Z(N111) );
  CKMUX2V8_8TH40 U15 ( .I0(n837), .I1(n832), .S(raddr2[4]), .Z(N171) );
  CKMUX2V8_8TH40 U16 ( .I0(n847), .I1(n842), .S(raddr2[4]), .Z(N170) );
  CKMUX2V8_8TH40 U17 ( .I0(n857), .I1(n852), .S(raddr2[4]), .Z(N169) );
  CKMUX2V8_8TH40 U18 ( .I0(n867), .I1(n862), .S(raddr2[4]), .Z(N168) );
  CKMUX2V8_8TH40 U19 ( .I0(n877), .I1(n872), .S(raddr2[4]), .Z(N167) );
  CKMUX2V8_8TH40 U20 ( .I0(n887), .I1(n882), .S(raddr2[4]), .Z(N166) );
  CKMUX2V8_8TH40 U21 ( .I0(n897), .I1(n892), .S(raddr2[4]), .Z(N165) );
  CKMUX2V8_8TH40 U22 ( .I0(n907), .I1(n902), .S(raddr2[4]), .Z(N164) );
  CKMUX2V8_8TH40 U23 ( .I0(n917), .I1(n912), .S(raddr2[4]), .Z(N163) );
  CKMUX2V8_8TH40 U24 ( .I0(n927), .I1(n922), .S(raddr2[4]), .Z(N162) );
  CKMUX2V8_8TH40 U25 ( .I0(n937), .I1(n932), .S(raddr2[4]), .Z(N161) );
  CKMUX2V8_8TH40 U26 ( .I0(n947), .I1(n942), .S(raddr2[4]), .Z(N160) );
  CKMUX2V8_8TH40 U27 ( .I0(n957), .I1(n952), .S(raddr2[4]), .Z(N159) );
  CKMUX2V8_8TH40 U28 ( .I0(n967), .I1(n962), .S(raddr2[4]), .Z(N158) );
  CKMUX2V8_8TH40 U29 ( .I0(n977), .I1(n972), .S(raddr2[4]), .Z(N157) );
  CKMUX2V8_8TH40 U30 ( .I0(n987), .I1(n982), .S(raddr2[4]), .Z(N156) );
  CKMUX2V8_8TH40 U31 ( .I0(n101), .I1(n96), .S(raddr1[4]), .Z(N126) );
  CKMUX2V8_8TH40 U32 ( .I0(n111), .I1(n106), .S(raddr1[4]), .Z(N125) );
  CKMUX2V8_8TH40 U33 ( .I0(n537), .I1(n532), .S(raddr1[4]), .Z(N124) );
  CKMUX2V8_8TH40 U34 ( .I0(n547), .I1(n542), .S(raddr1[4]), .Z(N123) );
  CKMUX2V8_8TH40 U35 ( .I0(n557), .I1(n552), .S(raddr1[4]), .Z(N122) );
  CKMUX2V8_8TH40 U36 ( .I0(n997), .I1(n992), .S(raddr2[4]), .Z(N155) );
  CKMUX2V8_8TH40 U37 ( .I0(n1007), .I1(n1002), .S(raddr2[4]), .Z(N154) );
  CKMUX2V8_8TH40 U38 ( .I0(n1017), .I1(n1012), .S(raddr2[4]), .Z(N153) );
  CKMUX2V8_8TH40 U39 ( .I0(n1027), .I1(n1022), .S(raddr2[4]), .Z(N152) );
  CKMUX2V8_8TH40 U40 ( .I0(n1037), .I1(n1032), .S(raddr2[4]), .Z(N151) );
  CKMUX2V8_8TH40 U41 ( .I0(n1047), .I1(n1042), .S(raddr2[4]), .Z(N150) );
  CKMUX2V8_8TH40 U42 ( .I0(n1057), .I1(n1052), .S(raddr2[4]), .Z(N149) );
  CKMUX2V8_8TH40 U43 ( .I0(n1067), .I1(n1062), .S(raddr2[4]), .Z(N148) );
  CKMUX2V8_8TH40 U44 ( .I0(n1077), .I1(n1072), .S(raddr2[4]), .Z(N147) );
  CKMUX2V8_8TH40 U45 ( .I0(n1087), .I1(n1082), .S(raddr2[4]), .Z(N146) );
  CKMUX2V8_8TH40 U46 ( .I0(n1097), .I1(n1092), .S(raddr2[4]), .Z(N145) );
  CKMUX2V8_8TH40 U47 ( .I0(n1107), .I1(n1102), .S(raddr2[4]), .Z(N144) );
  CKMUX2V8_8TH40 U48 ( .I0(n1117), .I1(n1112), .S(raddr2[4]), .Z(N143) );
  CKMUX2V8_8TH40 U49 ( .I0(n1127), .I1(n1122), .S(raddr2[4]), .Z(N142) );
  CKMUX2V8_8TH40 U50 ( .I0(n1137), .I1(n1132), .S(raddr2[4]), .Z(N141) );
  CKMUX2V8_8TH40 U51 ( .I0(n1147), .I1(n1142), .S(raddr2[4]), .Z(N140) );
  IOA22V4_8TH40 U52 ( .B1(n1171), .B2(n1193), .A1(N107), .A2(n1194), .ZN(
        rdata1[19]) );
  IOA22V4_8TH40 U53 ( .B1(n1172), .B2(n1193), .A1(N108), .A2(n1194), .ZN(
        rdata1[18]) );
  IOA22V4_8TH40 U54 ( .B1(n1173), .B2(n1193), .A1(N109), .A2(n1194), .ZN(
        rdata1[17]) );
  IOA22V4_8TH40 U55 ( .B1(n1174), .B2(n1193), .A1(N110), .A2(n1194), .ZN(
        rdata1[16]) );
  IOA22V4_8TH40 U56 ( .B1(n1157), .B2(n1193), .A1(N95), .A2(n1194), .ZN(
        rdata1[31]) );
  IOA22V4_8TH40 U57 ( .B1(n1158), .B2(n1193), .A1(N96), .A2(n1194), .ZN(
        rdata1[30]) );
  IOA22V4_8TH40 U58 ( .B1(n1160), .B2(n1193), .A1(N97), .A2(n1194), .ZN(
        rdata1[29]) );
  IOA22V4_8TH40 U59 ( .B1(n1161), .B2(n1193), .A1(N98), .A2(n1194), .ZN(
        rdata1[28]) );
  IOA22V4_8TH40 U60 ( .B1(n1162), .B2(n1193), .A1(N99), .A2(n1194), .ZN(
        rdata1[27]) );
  IOA22V4_8TH40 U61 ( .B1(n1163), .B2(n1193), .A1(N100), .A2(n1194), .ZN(
        rdata1[26]) );
  IOA22V4_8TH40 U62 ( .B1(n1164), .B2(n1193), .A1(N101), .A2(n1194), .ZN(
        rdata1[25]) );
  IOA22V4_8TH40 U63 ( .B1(n1165), .B2(n1193), .A1(N102), .A2(n1194), .ZN(
        rdata1[24]) );
  IOA22V4_8TH40 U64 ( .B1(n1166), .B2(n1193), .A1(N103), .A2(n1194), .ZN(
        rdata1[23]) );
  IOA22V4_8TH40 U65 ( .B1(n1167), .B2(n1193), .A1(N104), .A2(n1194), .ZN(
        rdata1[22]) );
  IOA22V4_8TH40 U66 ( .B1(n1168), .B2(n1193), .A1(N105), .A2(n1194), .ZN(
        rdata1[21]) );
  IOA22V4_8TH40 U67 ( .B1(n1169), .B2(n1193), .A1(N106), .A2(n1194), .ZN(
        rdata1[20]) );
  INOR2V2_8TH40 U68 ( .A1(n1220), .B1(n1210), .ZN(n1228) );
  INOR2V2_8TH40 U69 ( .A1(n1213), .B1(n1214), .ZN(n1231) );
  INOR2V2_8TH40 U70 ( .A1(n1212), .B1(n1208), .ZN(n1225) );
  INOR2V2_8TH40 U71 ( .A1(n1211), .B1(n1205), .ZN(n1216) );
  INOR2V2_8TH40 U72 ( .A1(n1220), .B1(n1214), .ZN(n1232) );
  INOR2V2_8TH40 U73 ( .A1(n1211), .B1(n1208), .ZN(n1224) );
  INOR2V2_8TH40 U74 ( .A1(n1212), .B1(n1205), .ZN(n1217) );
  INOR2V2_8TH40 U75 ( .A1(n1211), .B1(n1214), .ZN(n1229) );
  INOR2V2_8TH40 U76 ( .A1(n1220), .B1(n1208), .ZN(n1227) );
  INOR2V2_8TH40 U77 ( .A1(n1213), .B1(n1205), .ZN(n1218) );
  INOR2V2_8TH40 U78 ( .A1(n1212), .B1(n1214), .ZN(n1230) );
  INOR2V2_8TH40 U79 ( .A1(n1213), .B1(n1208), .ZN(n1226) );
  INOR2V2_8TH40 U80 ( .A1(n1220), .B1(n1205), .ZN(n1219) );
  INOR4V1_8TH40 U81 ( .A1(n1184), .B1(n3), .B2(raddr2[1]), .B3(raddr2[2]), 
        .ZN(n1183) );
  NOR2V0_8TH40 U82 ( .A1(raddr2[4]), .A2(raddr2[3]), .ZN(n1184) );
  INOR2V2_8TH40 U83 ( .A1(n1213), .B1(n1210), .ZN(n1246) );
  INOR2V2_8TH40 U84 ( .A1(n1212), .B1(n1210), .ZN(n1245) );
  INOR2V2_8TH40 U85 ( .A1(n1211), .B1(n1210), .ZN(n1243) );
  NOR2V2_8TH40 U86 ( .A1(n1205), .A2(n1207), .ZN(n1235) );
  NOR2V2_8TH40 U87 ( .A1(n1205), .A2(n1206), .ZN(n1234) );
  NOR2V2_8TH40 U88 ( .A1(n1207), .A2(n1214), .ZN(n1250) );
  NOR2V2_8TH40 U89 ( .A1(n1206), .A2(n1214), .ZN(n1249) );
  NOR2V2_8TH40 U90 ( .A1(n1204), .A2(n1214), .ZN(n1248) );
  NOR2V2_8TH40 U91 ( .A1(n1207), .A2(n1210), .ZN(n1244) );
  NOR2V2_8TH40 U92 ( .A1(n1206), .A2(n1210), .ZN(n1242) );
  NOR2V2_8TH40 U93 ( .A1(n1204), .A2(n1210), .ZN(n1241) );
  NOR2V2_8TH40 U94 ( .A1(n1207), .A2(n1208), .ZN(n1239) );
  NOR2V2_8TH40 U95 ( .A1(n1206), .A2(n1208), .ZN(n1238) );
  NOR2V2_8TH40 U96 ( .A1(n1204), .A2(n1208), .ZN(n1237) );
  NOR2V2_8TH40 U97 ( .A1(n1204), .A2(n1205), .ZN(n1233) );
  NOR2V2_8TH40 U98 ( .A1(n1209), .A2(n1214), .ZN(n1247) );
  NOR2V2_8TH40 U99 ( .A1(n1209), .A2(n1210), .ZN(n1240) );
  NOR2V2_8TH40 U100 ( .A1(n1208), .A2(n1209), .ZN(n1236) );
  NOR2V0_8TH40 U101 ( .A1(raddr1[4]), .A2(raddr1[3]), .ZN(n1197) );
  MOAI22V2_8TH40 U102 ( .A1(n1148), .A2(n1181), .B1(N171), .B2(n1150), .ZN(
        rdata2[0]) );
  MOAI22V2_8TH40 U103 ( .A1(n1148), .A2(n1170), .B1(N170), .B2(n1150), .ZN(
        rdata2[1]) );
  MOAI22V2_8TH40 U104 ( .A1(n1148), .A2(n1159), .B1(N169), .B2(n1150), .ZN(
        rdata2[2]) );
  MOAI22V2_8TH40 U105 ( .A1(n1148), .A2(n1156), .B1(N168), .B2(n1150), .ZN(
        rdata2[3]) );
  MOAI22V2_8TH40 U106 ( .A1(n1148), .A2(n1155), .B1(N167), .B2(n1150), .ZN(
        rdata2[4]) );
  MOAI22V2_8TH40 U107 ( .A1(n1148), .A2(n1154), .B1(N166), .B2(n1150), .ZN(
        rdata2[5]) );
  MOAI22V2_8TH40 U108 ( .A1(n1148), .A2(n1153), .B1(N165), .B2(n1150), .ZN(
        rdata2[6]) );
  MOAI22V2_8TH40 U109 ( .A1(n1148), .A2(n1152), .B1(N164), .B2(n1150), .ZN(
        rdata2[7]) );
  MOAI22V2_8TH40 U110 ( .A1(n1148), .A2(n1151), .B1(N163), .B2(n1150), .ZN(
        rdata2[8]) );
  MOAI22V2_8TH40 U111 ( .A1(n1148), .A2(n1149), .B1(N162), .B2(n1150), .ZN(
        rdata2[9]) );
  MOAI22V2_8TH40 U112 ( .A1(n1148), .A2(n1180), .B1(N161), .B2(n1150), .ZN(
        rdata2[10]) );
  MOAI22V2_8TH40 U113 ( .A1(n1148), .A2(n1179), .B1(N160), .B2(n1150), .ZN(
        rdata2[11]) );
  MOAI22V2_8TH40 U114 ( .A1(n1148), .A2(n1178), .B1(N159), .B2(n1150), .ZN(
        rdata2[12]) );
  MOAI22V2_8TH40 U115 ( .A1(n1148), .A2(n1177), .B1(N158), .B2(n1150), .ZN(
        rdata2[13]) );
  MOAI22V2_8TH40 U116 ( .A1(n1148), .A2(n1176), .B1(N157), .B2(n1150), .ZN(
        rdata2[14]) );
  MOAI22V2_8TH40 U117 ( .A1(n1148), .A2(n1175), .B1(N156), .B2(n1150), .ZN(
        rdata2[15]) );
  MOAI22V2_8TH40 U118 ( .A1(n1153), .A2(n1193), .B1(N120), .B2(n1194), .ZN(
        rdata1[6]) );
  MOAI22V2_8TH40 U119 ( .A1(n1152), .A2(n1193), .B1(N119), .B2(n1194), .ZN(
        rdata1[7]) );
  MOAI22V2_8TH40 U120 ( .A1(n1151), .A2(n1193), .B1(N118), .B2(n1194), .ZN(
        rdata1[8]) );
  MOAI22V2_8TH40 U121 ( .A1(n1149), .A2(n1193), .B1(N117), .B2(n1194), .ZN(
        rdata1[9]) );
  MOAI22V2_8TH40 U122 ( .A1(n1180), .A2(n1193), .B1(N116), .B2(n1194), .ZN(
        rdata1[10]) );
  MOAI22V2_8TH40 U123 ( .A1(n1179), .A2(n1193), .B1(N115), .B2(n1194), .ZN(
        rdata1[11]) );
  MOAI22V2_8TH40 U124 ( .A1(n1178), .A2(n1193), .B1(N114), .B2(n1194), .ZN(
        rdata1[12]) );
  MOAI22V2_8TH40 U125 ( .A1(n1177), .A2(n1193), .B1(N113), .B2(n1194), .ZN(
        rdata1[13]) );
  MOAI22V2_8TH40 U126 ( .A1(n1176), .A2(n1193), .B1(N112), .B2(n1194), .ZN(
        rdata1[14]) );
  MOAI22V2_8TH40 U127 ( .A1(n1175), .A2(n1193), .B1(N111), .B2(n1194), .ZN(
        rdata1[15]) );
  I2NOR4V2_8TH40 U128 ( .A1(re2), .A2(we), .B1(n1189), .B2(n1190), .ZN(n1188)
         );
  NAND4V2_8TH40 U129 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(
        n1195) );
  I2NOR4V2_8TH40 U130 ( .A1(we), .A2(re1), .B1(n1202), .B2(n1203), .ZN(n1201)
         );
  NAND4V2_8TH40 U131 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(
        n1182) );
  INV2_8TH40 U132 ( .I(n21), .ZN(n1) );
  INV2_8TH40 U133 ( .I(n21), .ZN(n2) );
  INV2_8TH40 U134 ( .I(n20), .ZN(n3) );
  INV2_8TH40 U135 ( .I(n20), .ZN(n4) );
  INV2_8TH40 U136 ( .I(n19), .ZN(n5) );
  INV2_8TH40 U137 ( .I(n19), .ZN(n6) );
  INV2_8TH40 U138 ( .I(n18), .ZN(n7) );
  INV2_8TH40 U139 ( .I(n18), .ZN(n8) );
  INV2_8TH40 U140 ( .I(n17), .ZN(n9) );
  INV2_8TH40 U141 ( .I(n17), .ZN(n10) );
  INV2_8TH40 U142 ( .I(n16), .ZN(n11) );
  INV2_8TH40 U143 ( .I(n16), .ZN(n12) );
  INV2_8TH40 U144 ( .I(n15), .ZN(n13) );
  INV2_8TH40 U145 ( .I(n15), .ZN(n14) );
  INV2_8TH40 U146 ( .I(n66), .ZN(n45) );
  INV2_8TH40 U147 ( .I(n66), .ZN(n46) );
  INV2_8TH40 U148 ( .I(n65), .ZN(n47) );
  INV2_8TH40 U149 ( .I(n65), .ZN(n48) );
  INV2_8TH40 U150 ( .I(n64), .ZN(n49) );
  INV2_8TH40 U151 ( .I(n64), .ZN(n50) );
  INV2_8TH40 U152 ( .I(n63), .ZN(n51) );
  INV2_8TH40 U153 ( .I(n63), .ZN(n52) );
  INV2_8TH40 U154 ( .I(n62), .ZN(n53) );
  INV2_8TH40 U155 ( .I(n61), .ZN(n54) );
  INV2_8TH40 U156 ( .I(n60), .ZN(n55) );
  INV2_8TH40 U157 ( .I(n60), .ZN(n56) );
  INV2_8TH40 U158 ( .I(n59), .ZN(n57) );
  INV2_8TH40 U159 ( .I(n59), .ZN(n58) );
  INV2_8TH40 U160 ( .I(n39), .ZN(n31) );
  INV2_8TH40 U161 ( .I(n39), .ZN(n32) );
  INV2_8TH40 U162 ( .I(n38), .ZN(n33) );
  INV2_8TH40 U163 ( .I(n38), .ZN(n34) );
  INV2_8TH40 U164 ( .I(n37), .ZN(n35) );
  INV2_8TH40 U165 ( .I(n37), .ZN(n36) );
  INV2_8TH40 U166 ( .I(n43), .ZN(n23) );
  INV2_8TH40 U167 ( .I(n43), .ZN(n24) );
  INV2_8TH40 U168 ( .I(n42), .ZN(n25) );
  INV2_8TH40 U169 ( .I(n42), .ZN(n26) );
  INV2_8TH40 U170 ( .I(n41), .ZN(n27) );
  INV2_8TH40 U171 ( .I(n41), .ZN(n28) );
  INV2_8TH40 U172 ( .I(n40), .ZN(n29) );
  INV2_8TH40 U173 ( .I(n40), .ZN(n30) );
  CLKBUFV2_8TH40 U174 ( .I(n22), .Z(n21) );
  CLKBUFV2_8TH40 U175 ( .I(n22), .Z(n20) );
  CLKBUFV2_8TH40 U176 ( .I(n44), .Z(n39) );
  CLKBUFV2_8TH40 U177 ( .I(n17), .Z(n19) );
  CLKBUFV2_8TH40 U178 ( .I(n44), .Z(n38) );
  CLKBUFV2_8TH40 U179 ( .I(n16), .Z(n18) );
  CLKBUFV2_8TH40 U180 ( .I(n44), .Z(n37) );
  CLKBUFV2_8TH40 U181 ( .I(n21), .Z(n17) );
  CLKBUFV2_8TH40 U182 ( .I(n20), .Z(n16) );
  CLKBUFV2_8TH40 U183 ( .I(n41), .Z(n43) );
  CLKBUFV2_8TH40 U184 ( .I(n40), .Z(n42) );
  CLKBUFV2_8TH40 U185 ( .I(n39), .Z(n41) );
  CLKBUFV2_8TH40 U186 ( .I(n38), .Z(n40) );
  CLKBUFV2_8TH40 U187 ( .I(n22), .Z(n15) );
  CLKBUFV2_8TH40 U188 ( .I(n67), .Z(n66) );
  CLKBUFV2_8TH40 U189 ( .I(n67), .Z(n65) );
  CLKBUFV2_8TH40 U190 ( .I(n63), .Z(n64) );
  CLKBUFV2_8TH40 U191 ( .I(n66), .Z(n63) );
  CLKBUFV2_8TH40 U192 ( .I(n65), .Z(n62) );
  CLKBUFV2_8TH40 U193 ( .I(n60), .Z(n61) );
  CLKBUFV2_8TH40 U194 ( .I(n59), .Z(n60) );
  CLKBUFV2_8TH40 U195 ( .I(n67), .Z(n59) );
  INV2_8TH40 U196 ( .I(n87), .ZN(n74) );
  INV2_8TH40 U197 ( .I(n87), .ZN(n75) );
  INV2_8TH40 U198 ( .I(n86), .ZN(n76) );
  INV2_8TH40 U199 ( .I(n86), .ZN(n77) );
  INV2_8TH40 U200 ( .I(n85), .ZN(n78) );
  INV2_8TH40 U201 ( .I(n85), .ZN(n79) );
  INV2_8TH40 U202 ( .I(n84), .ZN(n80) );
  INV2_8TH40 U203 ( .I(n84), .ZN(n81) );
  INV2_8TH40 U204 ( .I(n83), .ZN(n82) );
  INV2_8TH40 U205 ( .I(n90), .ZN(n68) );
  INV2_8TH40 U206 ( .I(n90), .ZN(n69) );
  INV2_8TH40 U207 ( .I(n89), .ZN(n70) );
  INV2_8TH40 U208 ( .I(n89), .ZN(n71) );
  INV2_8TH40 U209 ( .I(n88), .ZN(n72) );
  INV2_8TH40 U210 ( .I(n88), .ZN(n73) );
  INV2_8TH40 U211 ( .I(raddr2[0]), .ZN(n22) );
  INV2_8TH40 U212 ( .I(raddr2[1]), .ZN(n44) );
  INV2_8TH40 U213 ( .I(raddr1[0]), .ZN(n67) );
  CLKBUFV2_8TH40 U214 ( .I(n86), .Z(n87) );
  CLKBUFV2_8TH40 U215 ( .I(n91), .Z(n86) );
  CLKBUFV2_8TH40 U216 ( .I(n91), .Z(n85) );
  CLKBUFV2_8TH40 U217 ( .I(n83), .Z(n84) );
  CLKBUFV2_8TH40 U218 ( .I(n91), .Z(n83) );
  CLKBUFV2_8TH40 U219 ( .I(n87), .Z(n90) );
  CLKBUFV2_8TH40 U220 ( .I(n88), .Z(n89) );
  CLKBUFV2_8TH40 U221 ( .I(n85), .Z(n88) );
  INV2_8TH40 U222 ( .I(raddr1[1]), .ZN(n91) );
  MUX4V2_8TH40 U223 ( .I0(regs[624]), .I1(regs[592]), .I2(regs[560]), .I3(
        regs[528]), .S0(n53), .S1(n68), .Z(n673) );
  MUX4V2_8TH40 U224 ( .I0(regs[880]), .I1(regs[848]), .I2(regs[816]), .I3(
        regs[784]), .S0(n53), .S1(n68), .Z(n675) );
  MUX4V2_8TH40 U225 ( .I0(regs[1008]), .I1(regs[976]), .I2(regs[944]), .I3(
        regs[912]), .S0(n53), .S1(n68), .Z(n676) );
  MUX4V2_8TH40 U226 ( .I0(regs[625]), .I1(regs[593]), .I2(regs[561]), .I3(
        regs[529]), .S0(n53), .S1(n68), .Z(n683) );
  MUX4V2_8TH40 U227 ( .I0(regs[881]), .I1(regs[849]), .I2(regs[817]), .I3(
        regs[785]), .S0(n53), .S1(n69), .Z(n685) );
  MUX4V2_8TH40 U228 ( .I0(regs[1009]), .I1(regs[977]), .I2(regs[945]), .I3(
        regs[913]), .S0(n58), .S1(n69), .Z(n686) );
  MUX4V2_8TH40 U229 ( .I0(regs[626]), .I1(regs[594]), .I2(regs[562]), .I3(
        regs[530]), .S0(n51), .S1(n69), .Z(n693) );
  MUX4V2_8TH40 U230 ( .I0(regs[882]), .I1(regs[850]), .I2(regs[818]), .I3(
        regs[786]), .S0(n50), .S1(n69), .Z(n695) );
  MUX4V2_8TH40 U231 ( .I0(regs[1010]), .I1(regs[978]), .I2(regs[946]), .I3(
        regs[914]), .S0(n49), .S1(n69), .Z(n696) );
  MUX4V2_8TH40 U232 ( .I0(regs[627]), .I1(regs[595]), .I2(regs[563]), .I3(
        regs[531]), .S0(n54), .S1(n70), .Z(n703) );
  MUX4V2_8TH40 U233 ( .I0(regs[883]), .I1(regs[851]), .I2(regs[819]), .I3(
        regs[787]), .S0(n54), .S1(n70), .Z(n705) );
  MUX4V2_8TH40 U234 ( .I0(regs[1011]), .I1(regs[979]), .I2(regs[947]), .I3(
        regs[915]), .S0(n54), .S1(n70), .Z(n706) );
  MUX4V2_8TH40 U235 ( .I0(regs[628]), .I1(regs[596]), .I2(regs[564]), .I3(
        regs[532]), .S0(n54), .S1(n70), .Z(n713) );
  MUX4V2_8TH40 U236 ( .I0(regs[884]), .I1(regs[852]), .I2(regs[820]), .I3(
        regs[788]), .S0(n54), .S1(n70), .Z(n715) );
  MUX4V2_8TH40 U237 ( .I0(regs[1012]), .I1(regs[980]), .I2(regs[948]), .I3(
        regs[916]), .S0(n54), .S1(n71), .Z(n716) );
  MUX4V2_8TH40 U238 ( .I0(regs[629]), .I1(regs[597]), .I2(regs[565]), .I3(
        regs[533]), .S0(n57), .S1(n71), .Z(n723) );
  MUX4V2_8TH40 U239 ( .I0(regs[885]), .I1(regs[853]), .I2(regs[821]), .I3(
        regs[789]), .S0(n48), .S1(n71), .Z(n725) );
  MUX4V2_8TH40 U240 ( .I0(regs[1013]), .I1(regs[981]), .I2(regs[949]), .I3(
        regs[917]), .S0(n47), .S1(n71), .Z(n726) );
  MUX4V2_8TH40 U241 ( .I0(regs[630]), .I1(regs[598]), .I2(regs[566]), .I3(
        regs[534]), .S0(n58), .S1(n81), .Z(n733) );
  MUX4V2_8TH40 U242 ( .I0(regs[886]), .I1(regs[854]), .I2(regs[822]), .I3(
        regs[790]), .S0(n55), .S1(n80), .Z(n735) );
  MUX4V2_8TH40 U243 ( .I0(regs[1014]), .I1(regs[982]), .I2(regs[950]), .I3(
        regs[918]), .S0(n55), .S1(n82), .Z(n736) );
  MUX4V2_8TH40 U244 ( .I0(regs[631]), .I1(regs[599]), .I2(regs[567]), .I3(
        regs[535]), .S0(n55), .S1(raddr1[1]), .Z(n743) );
  MUX4V2_8TH40 U245 ( .I0(regs[887]), .I1(regs[855]), .I2(regs[823]), .I3(
        regs[791]), .S0(n55), .S1(n71), .Z(n745) );
  MUX4V2_8TH40 U246 ( .I0(regs[1015]), .I1(regs[983]), .I2(regs[951]), .I3(
        regs[919]), .S0(n55), .S1(n77), .Z(n746) );
  MUX4V2_8TH40 U247 ( .I0(regs[632]), .I1(regs[600]), .I2(regs[568]), .I3(
        regs[536]), .S0(n56), .S1(n69), .Z(n753) );
  MUX4V2_8TH40 U248 ( .I0(regs[888]), .I1(regs[856]), .I2(regs[824]), .I3(
        regs[792]), .S0(n56), .S1(n68), .Z(n755) );
  MUX4V2_8TH40 U249 ( .I0(regs[1016]), .I1(regs[984]), .I2(regs[952]), .I3(
        regs[920]), .S0(n56), .S1(raddr1[1]), .Z(n756) );
  MUX4V2_8TH40 U250 ( .I0(regs[633]), .I1(regs[601]), .I2(regs[569]), .I3(
        regs[537]), .S0(n56), .S1(n74), .Z(n763) );
  MUX4V2_8TH40 U251 ( .I0(regs[889]), .I1(regs[857]), .I2(regs[825]), .I3(
        regs[793]), .S0(n56), .S1(n71), .Z(n765) );
  MUX4V2_8TH40 U252 ( .I0(regs[1017]), .I1(regs[985]), .I2(regs[953]), .I3(
        regs[921]), .S0(n56), .S1(n70), .Z(n766) );
  MUX4V2_8TH40 U253 ( .I0(regs[634]), .I1(regs[602]), .I2(regs[570]), .I3(
        regs[538]), .S0(n57), .S1(n78), .Z(n773) );
  MUX4V2_8TH40 U254 ( .I0(regs[890]), .I1(regs[858]), .I2(regs[826]), .I3(
        regs[794]), .S0(n57), .S1(n73), .Z(n775) );
  MUX4V2_8TH40 U255 ( .I0(regs[1018]), .I1(regs[986]), .I2(regs[954]), .I3(
        regs[922]), .S0(n57), .S1(n72), .Z(n776) );
  MUX4V2_8TH40 U256 ( .I0(regs[635]), .I1(regs[603]), .I2(regs[571]), .I3(
        regs[539]), .S0(n57), .S1(n78), .Z(n783) );
  MUX4V2_8TH40 U257 ( .I0(regs[891]), .I1(regs[859]), .I2(regs[827]), .I3(
        regs[795]), .S0(n58), .S1(n73), .Z(n785) );
  MUX4V2_8TH40 U258 ( .I0(regs[1019]), .I1(regs[987]), .I2(regs[955]), .I3(
        regs[923]), .S0(n58), .S1(n72), .Z(n786) );
  MUX4V2_8TH40 U259 ( .I0(regs[636]), .I1(regs[604]), .I2(regs[572]), .I3(
        regs[540]), .S0(n58), .S1(n80), .Z(n793) );
  MUX4V2_8TH40 U260 ( .I0(regs[892]), .I1(regs[860]), .I2(regs[828]), .I3(
        regs[796]), .S0(n58), .S1(n82), .Z(n795) );
  MUX4V2_8TH40 U261 ( .I0(regs[1020]), .I1(regs[988]), .I2(regs[956]), .I3(
        regs[924]), .S0(n58), .S1(n79), .Z(n796) );
  MUX4V2_8TH40 U262 ( .I0(regs[637]), .I1(regs[605]), .I2(regs[573]), .I3(
        regs[541]), .S0(raddr1[0]), .S1(n72), .Z(n803) );
  MUX4V2_8TH40 U263 ( .I0(regs[893]), .I1(regs[861]), .I2(regs[829]), .I3(
        regs[797]), .S0(raddr1[0]), .S1(n72), .Z(n805) );
  MUX4V2_8TH40 U264 ( .I0(regs[1021]), .I1(regs[989]), .I2(regs[957]), .I3(
        regs[925]), .S0(raddr1[0]), .S1(n72), .Z(n806) );
  MUX4V2_8TH40 U265 ( .I0(regs[638]), .I1(regs[606]), .I2(regs[574]), .I3(
        regs[542]), .S0(n50), .S1(n72), .Z(n813) );
  MUX4V2_8TH40 U266 ( .I0(regs[894]), .I1(regs[862]), .I2(regs[830]), .I3(
        regs[798]), .S0(n49), .S1(n73), .Z(n815) );
  MUX4V2_8TH40 U267 ( .I0(regs[1022]), .I1(regs[990]), .I2(regs[958]), .I3(
        regs[926]), .S0(raddr1[0]), .S1(n73), .Z(n816) );
  MUX4V2_8TH40 U268 ( .I0(regs[639]), .I1(regs[607]), .I2(regs[575]), .I3(
        regs[543]), .S0(raddr1[0]), .S1(n73), .Z(n823) );
  MUX4V2_8TH40 U269 ( .I0(regs[895]), .I1(regs[863]), .I2(regs[831]), .I3(
        regs[799]), .S0(raddr1[0]), .S1(n73), .Z(n825) );
  MUX4V2_8TH40 U270 ( .I0(regs[1023]), .I1(regs[991]), .I2(regs[959]), .I3(
        regs[927]), .S0(raddr1[0]), .S1(n73), .Z(n826) );
  MUX4V2_8TH40 U271 ( .I0(regs[101]), .I1(regs[69]), .I2(regs[37]), .I3(
        regs[5]), .S0(n48), .S1(n76), .Z(n558) );
  MUX4V2_8TH40 U272 ( .I0(regs[102]), .I1(regs[70]), .I2(regs[38]), .I3(
        regs[6]), .S0(n48), .S1(n77), .Z(n568) );
  MUX4V2_8TH40 U273 ( .I0(regs[103]), .I1(regs[71]), .I2(regs[39]), .I3(
        regs[7]), .S0(n49), .S1(n78), .Z(n578) );
  MUX4V2_8TH40 U274 ( .I0(regs[104]), .I1(regs[72]), .I2(regs[40]), .I3(
        regs[8]), .S0(n49), .S1(n78), .Z(n588) );
  MUX4V2_8TH40 U275 ( .I0(regs[105]), .I1(regs[73]), .I2(regs[41]), .I3(
        regs[9]), .S0(n50), .S1(n79), .Z(n598) );
  MUX4V2_8TH40 U276 ( .I0(regs[106]), .I1(regs[74]), .I2(regs[42]), .I3(
        regs[10]), .S0(n58), .S1(n79), .Z(n608) );
  MUX4V2_8TH40 U277 ( .I0(regs[107]), .I1(regs[75]), .I2(regs[43]), .I3(
        regs[11]), .S0(n49), .S1(n80), .Z(n618) );
  MUX4V2_8TH40 U278 ( .I0(regs[108]), .I1(regs[76]), .I2(regs[44]), .I3(
        regs[12]), .S0(n55), .S1(n81), .Z(n628) );
  MUX4V2_8TH40 U279 ( .I0(regs[109]), .I1(regs[77]), .I2(regs[45]), .I3(
        regs[13]), .S0(n51), .S1(n81), .Z(n638) );
  MUX4V2_8TH40 U280 ( .I0(regs[110]), .I1(regs[78]), .I2(regs[46]), .I3(
        regs[14]), .S0(n51), .S1(n82), .Z(n648) );
  MUX4V2_8TH40 U281 ( .I0(regs[111]), .I1(regs[79]), .I2(regs[47]), .I3(
        regs[15]), .S0(n52), .S1(raddr1[1]), .Z(n658) );
  MUX4V2_8TH40 U282 ( .I0(regs[96]), .I1(regs[64]), .I2(regs[32]), .I3(regs[0]), .S0(n1), .S1(n23), .Z(n828) );
  MUX4V2_8TH40 U283 ( .I0(regs[97]), .I1(regs[65]), .I2(regs[33]), .I3(regs[1]), .S0(n1), .S1(n29), .Z(n838) );
  MUX4V2_8TH40 U284 ( .I0(regs[98]), .I1(regs[66]), .I2(regs[34]), .I3(regs[2]), .S0(n2), .S1(n35), .Z(n848) );
  MUX4V2_8TH40 U285 ( .I0(regs[99]), .I1(regs[67]), .I2(regs[35]), .I3(regs[3]), .S0(n2), .S1(n36), .Z(n858) );
  MUX4V2_8TH40 U286 ( .I0(regs[100]), .I1(regs[68]), .I2(regs[36]), .I3(
        regs[4]), .S0(n3), .S1(n31), .Z(n868) );
  MUX4V2_8TH40 U287 ( .I0(regs[101]), .I1(regs[69]), .I2(regs[37]), .I3(
        regs[5]), .S0(n4), .S1(n31), .Z(n878) );
  MUX4V2_8TH40 U288 ( .I0(regs[102]), .I1(regs[70]), .I2(regs[38]), .I3(
        regs[6]), .S0(n4), .S1(n32), .Z(n888) );
  MUX4V2_8TH40 U289 ( .I0(regs[103]), .I1(regs[71]), .I2(regs[39]), .I3(
        regs[7]), .S0(n5), .S1(n33), .Z(n898) );
  MUX4V2_8TH40 U290 ( .I0(regs[104]), .I1(regs[72]), .I2(regs[40]), .I3(
        regs[8]), .S0(n5), .S1(n33), .Z(n908) );
  MUX4V2_8TH40 U291 ( .I0(regs[105]), .I1(regs[73]), .I2(regs[41]), .I3(
        regs[9]), .S0(n6), .S1(n34), .Z(n918) );
  MUX4V2_8TH40 U292 ( .I0(regs[106]), .I1(regs[74]), .I2(regs[42]), .I3(
        regs[10]), .S0(n7), .S1(n34), .Z(n928) );
  MUX4V2_8TH40 U293 ( .I0(regs[107]), .I1(regs[75]), .I2(regs[43]), .I3(
        regs[11]), .S0(n7), .S1(n35), .Z(n938) );
  MUX4V2_8TH40 U294 ( .I0(regs[108]), .I1(regs[76]), .I2(regs[44]), .I3(
        regs[12]), .S0(n8), .S1(n36), .Z(n948) );
  MUX4V2_8TH40 U295 ( .I0(regs[109]), .I1(regs[77]), .I2(regs[45]), .I3(
        regs[13]), .S0(n9), .S1(n36), .Z(n958) );
  MUX4V2_8TH40 U296 ( .I0(regs[110]), .I1(regs[78]), .I2(regs[46]), .I3(
        regs[14]), .S0(n9), .S1(raddr2[1]), .Z(n968) );
  MUX4V2_8TH40 U297 ( .I0(regs[111]), .I1(regs[79]), .I2(regs[47]), .I3(
        regs[15]), .S0(n10), .S1(raddr2[1]), .Z(n978) );
  MUX4V2_8TH40 U298 ( .I0(regs[736]), .I1(regs[704]), .I2(regs[672]), .I3(
        regs[640]), .S0(n1), .S1(n30), .Z(n834) );
  MUX4V2_8TH40 U299 ( .I0(regs[224]), .I1(regs[192]), .I2(regs[160]), .I3(
        regs[128]), .S0(n1), .S1(n33), .Z(n829) );
  MUX4V2_8TH40 U300 ( .I0(regs[737]), .I1(regs[705]), .I2(regs[673]), .I3(
        regs[641]), .S0(n2), .S1(n33), .Z(n844) );
  MUX4V2_8TH40 U301 ( .I0(regs[225]), .I1(regs[193]), .I2(regs[161]), .I3(
        regs[129]), .S0(n1), .S1(n34), .Z(n839) );
  MUX4V2_8TH40 U302 ( .I0(regs[738]), .I1(regs[706]), .I2(regs[674]), .I3(
        regs[642]), .S0(n2), .S1(n32), .Z(n854) );
  MUX4V2_8TH40 U303 ( .I0(regs[226]), .I1(regs[194]), .I2(regs[162]), .I3(
        regs[130]), .S0(n2), .S1(n32), .Z(n849) );
  MUX4V2_8TH40 U304 ( .I0(regs[739]), .I1(regs[707]), .I2(regs[675]), .I3(
        regs[643]), .S0(n3), .S1(n31), .Z(n864) );
  MUX4V2_8TH40 U305 ( .I0(regs[227]), .I1(regs[195]), .I2(regs[163]), .I3(
        regs[131]), .S0(n2), .S1(n26), .Z(n859) );
  MUX4V2_8TH40 U306 ( .I0(regs[740]), .I1(regs[708]), .I2(regs[676]), .I3(
        regs[644]), .S0(n3), .S1(n31), .Z(n874) );
  MUX4V2_8TH40 U307 ( .I0(regs[228]), .I1(regs[196]), .I2(regs[164]), .I3(
        regs[132]), .S0(n3), .S1(n31), .Z(n869) );
  MUX4V2_8TH40 U308 ( .I0(regs[741]), .I1(regs[709]), .I2(regs[677]), .I3(
        regs[645]), .S0(n4), .S1(n32), .Z(n884) );
  MUX4V2_8TH40 U309 ( .I0(regs[229]), .I1(regs[197]), .I2(regs[165]), .I3(
        regs[133]), .S0(n4), .S1(n31), .Z(n879) );
  MUX4V2_8TH40 U310 ( .I0(regs[742]), .I1(regs[710]), .I2(regs[678]), .I3(
        regs[646]), .S0(n5), .S1(n32), .Z(n894) );
  MUX4V2_8TH40 U311 ( .I0(regs[230]), .I1(regs[198]), .I2(regs[166]), .I3(
        regs[134]), .S0(n4), .S1(n32), .Z(n889) );
  MUX4V2_8TH40 U312 ( .I0(regs[743]), .I1(regs[711]), .I2(regs[679]), .I3(
        regs[647]), .S0(n5), .S1(n33), .Z(n904) );
  MUX4V2_8TH40 U313 ( .I0(regs[231]), .I1(regs[199]), .I2(regs[167]), .I3(
        regs[135]), .S0(n5), .S1(n33), .Z(n899) );
  MUX4V2_8TH40 U314 ( .I0(regs[744]), .I1(regs[712]), .I2(regs[680]), .I3(
        regs[648]), .S0(n6), .S1(n34), .Z(n914) );
  MUX4V2_8TH40 U315 ( .I0(regs[232]), .I1(regs[200]), .I2(regs[168]), .I3(
        regs[136]), .S0(n6), .S1(n33), .Z(n909) );
  MUX4V2_8TH40 U316 ( .I0(regs[745]), .I1(regs[713]), .I2(regs[681]), .I3(
        regs[649]), .S0(n6), .S1(n34), .Z(n924) );
  MUX4V2_8TH40 U317 ( .I0(regs[233]), .I1(regs[201]), .I2(regs[169]), .I3(
        regs[137]), .S0(n6), .S1(n34), .Z(n919) );
  MUX4V2_8TH40 U318 ( .I0(regs[746]), .I1(regs[714]), .I2(regs[682]), .I3(
        regs[650]), .S0(n7), .S1(n35), .Z(n934) );
  MUX4V2_8TH40 U319 ( .I0(regs[234]), .I1(regs[202]), .I2(regs[170]), .I3(
        regs[138]), .S0(n7), .S1(n35), .Z(n929) );
  MUX4V2_8TH40 U320 ( .I0(regs[747]), .I1(regs[715]), .I2(regs[683]), .I3(
        regs[651]), .S0(n8), .S1(n36), .Z(n944) );
  MUX4V2_8TH40 U321 ( .I0(regs[235]), .I1(regs[203]), .I2(regs[171]), .I3(
        regs[139]), .S0(n7), .S1(n35), .Z(n939) );
  MUX4V2_8TH40 U322 ( .I0(regs[748]), .I1(regs[716]), .I2(regs[684]), .I3(
        regs[652]), .S0(n8), .S1(n36), .Z(n954) );
  MUX4V2_8TH40 U323 ( .I0(regs[236]), .I1(regs[204]), .I2(regs[172]), .I3(
        regs[140]), .S0(n8), .S1(n36), .Z(n949) );
  MUX4V2_8TH40 U324 ( .I0(regs[749]), .I1(regs[717]), .I2(regs[685]), .I3(
        regs[653]), .S0(n9), .S1(n23), .Z(n964) );
  MUX4V2_8TH40 U325 ( .I0(regs[237]), .I1(regs[205]), .I2(regs[173]), .I3(
        regs[141]), .S0(n9), .S1(n24), .Z(n959) );
  MUX4V2_8TH40 U326 ( .I0(regs[750]), .I1(regs[718]), .I2(regs[686]), .I3(
        regs[654]), .S0(n10), .S1(n27), .Z(n974) );
  MUX4V2_8TH40 U327 ( .I0(regs[238]), .I1(regs[206]), .I2(regs[174]), .I3(
        regs[142]), .S0(n9), .S1(n28), .Z(n969) );
  MUX4V2_8TH40 U328 ( .I0(regs[751]), .I1(regs[719]), .I2(regs[687]), .I3(
        regs[655]), .S0(n10), .S1(raddr2[1]), .Z(n984) );
  MUX4V2_8TH40 U329 ( .I0(regs[239]), .I1(regs[207]), .I2(regs[175]), .I3(
        regs[143]), .S0(n10), .S1(raddr2[1]), .Z(n979) );
  MUX4V2_8TH40 U330 ( .I0(regs[752]), .I1(regs[720]), .I2(regs[688]), .I3(
        regs[656]), .S0(n11), .S1(n23), .Z(n994) );
  MUX4V2_8TH40 U331 ( .I0(regs[240]), .I1(regs[208]), .I2(regs[176]), .I3(
        regs[144]), .S0(n10), .S1(n23), .Z(n989) );
  MUX4V2_8TH40 U332 ( .I0(regs[753]), .I1(regs[721]), .I2(regs[689]), .I3(
        regs[657]), .S0(n11), .S1(n24), .Z(n1004) );
  MUX4V2_8TH40 U333 ( .I0(regs[241]), .I1(regs[209]), .I2(regs[177]), .I3(
        regs[145]), .S0(n11), .S1(n23), .Z(n999) );
  MUX4V2_8TH40 U334 ( .I0(regs[754]), .I1(regs[722]), .I2(regs[690]), .I3(
        regs[658]), .S0(n12), .S1(n24), .Z(n1014) );
  MUX4V2_8TH40 U335 ( .I0(regs[242]), .I1(regs[210]), .I2(regs[178]), .I3(
        regs[146]), .S0(n12), .S1(n24), .Z(n1009) );
  MUX4V2_8TH40 U336 ( .I0(regs[755]), .I1(regs[723]), .I2(regs[691]), .I3(
        regs[659]), .S0(n7), .S1(n25), .Z(n1024) );
  MUX4V2_8TH40 U337 ( .I0(regs[243]), .I1(regs[211]), .I2(regs[179]), .I3(
        regs[147]), .S0(n12), .S1(n24), .Z(n1019) );
  MUX4V2_8TH40 U338 ( .I0(regs[756]), .I1(regs[724]), .I2(regs[692]), .I3(
        regs[660]), .S0(n8), .S1(n25), .Z(n1034) );
  MUX4V2_8TH40 U339 ( .I0(regs[244]), .I1(regs[212]), .I2(regs[180]), .I3(
        regs[148]), .S0(n11), .S1(n25), .Z(n1029) );
  MUX4V2_8TH40 U340 ( .I0(regs[757]), .I1(regs[725]), .I2(regs[693]), .I3(
        regs[661]), .S0(n13), .S1(n26), .Z(n1044) );
  MUX4V2_8TH40 U341 ( .I0(regs[245]), .I1(regs[213]), .I2(regs[181]), .I3(
        regs[149]), .S0(n14), .S1(n26), .Z(n1039) );
  MUX4V2_8TH40 U342 ( .I0(regs[758]), .I1(regs[726]), .I2(regs[694]), .I3(
        regs[662]), .S0(n10), .S1(n27), .Z(n1054) );
  MUX4V2_8TH40 U343 ( .I0(regs[246]), .I1(regs[214]), .I2(regs[182]), .I3(
        regs[150]), .S0(n10), .S1(n26), .Z(n1049) );
  MUX4V2_8TH40 U344 ( .I0(regs[759]), .I1(regs[727]), .I2(regs[695]), .I3(
        regs[663]), .S0(n1), .S1(n27), .Z(n1064) );
  MUX4V2_8TH40 U345 ( .I0(regs[247]), .I1(regs[215]), .I2(regs[183]), .I3(
        regs[151]), .S0(n2), .S1(n27), .Z(n1059) );
  MUX4V2_8TH40 U346 ( .I0(regs[760]), .I1(regs[728]), .I2(regs[696]), .I3(
        regs[664]), .S0(n1), .S1(n28), .Z(n1074) );
  MUX4V2_8TH40 U347 ( .I0(regs[248]), .I1(regs[216]), .I2(regs[184]), .I3(
        regs[152]), .S0(n7), .S1(n25), .Z(n1069) );
  MUX4V2_8TH40 U348 ( .I0(regs[761]), .I1(regs[729]), .I2(regs[697]), .I3(
        regs[665]), .S0(n2), .S1(n28), .Z(n1084) );
  MUX4V2_8TH40 U349 ( .I0(regs[249]), .I1(regs[217]), .I2(regs[185]), .I3(
        regs[153]), .S0(n7), .S1(n28), .Z(n1079) );
  MUX4V2_8TH40 U350 ( .I0(regs[762]), .I1(regs[730]), .I2(regs[698]), .I3(
        regs[666]), .S0(n13), .S1(n29), .Z(n1094) );
  MUX4V2_8TH40 U351 ( .I0(regs[250]), .I1(regs[218]), .I2(regs[186]), .I3(
        regs[154]), .S0(n13), .S1(n29), .Z(n1089) );
  MUX4V2_8TH40 U352 ( .I0(regs[763]), .I1(regs[731]), .I2(regs[699]), .I3(
        regs[667]), .S0(n14), .S1(n30), .Z(n1104) );
  MUX4V2_8TH40 U353 ( .I0(regs[251]), .I1(regs[219]), .I2(regs[187]), .I3(
        regs[155]), .S0(n13), .S1(n29), .Z(n1099) );
  MUX4V2_8TH40 U354 ( .I0(regs[764]), .I1(regs[732]), .I2(regs[700]), .I3(
        regs[668]), .S0(n14), .S1(n30), .Z(n1114) );
  MUX4V2_8TH40 U355 ( .I0(regs[252]), .I1(regs[220]), .I2(regs[188]), .I3(
        regs[156]), .S0(n14), .S1(n30), .Z(n1109) );
  MUX4V2_8TH40 U356 ( .I0(regs[765]), .I1(regs[733]), .I2(regs[701]), .I3(
        regs[669]), .S0(raddr2[0]), .S1(n25), .Z(n1124) );
  MUX4V2_8TH40 U357 ( .I0(regs[253]), .I1(regs[221]), .I2(regs[189]), .I3(
        regs[157]), .S0(n14), .S1(n26), .Z(n1119) );
  MUX4V2_8TH40 U358 ( .I0(regs[766]), .I1(regs[734]), .I2(regs[702]), .I3(
        regs[670]), .S0(raddr2[0]), .S1(n26), .Z(n1134) );
  MUX4V2_8TH40 U359 ( .I0(regs[254]), .I1(regs[222]), .I2(regs[190]), .I3(
        regs[158]), .S0(raddr2[0]), .S1(n29), .Z(n1129) );
  MUX4V2_8TH40 U360 ( .I0(regs[736]), .I1(regs[704]), .I2(regs[672]), .I3(
        regs[640]), .S0(n45), .S1(n74), .Z(n98) );
  MUX4V2_8TH40 U361 ( .I0(regs[224]), .I1(regs[192]), .I2(regs[160]), .I3(
        regs[128]), .S0(n45), .S1(n78), .Z(n93) );
  MUX4V2_8TH40 U362 ( .I0(regs[737]), .I1(regs[705]), .I2(regs[673]), .I3(
        regs[641]), .S0(n46), .S1(n74), .Z(n108) );
  MUX4V2_8TH40 U363 ( .I0(regs[225]), .I1(regs[193]), .I2(regs[161]), .I3(
        regs[129]), .S0(n45), .S1(n74), .Z(n103) );
  MUX4V2_8TH40 U364 ( .I0(regs[738]), .I1(regs[706]), .I2(regs[674]), .I3(
        regs[642]), .S0(n46), .S1(n75), .Z(n534) );
  MUX4V2_8TH40 U365 ( .I0(regs[226]), .I1(regs[194]), .I2(regs[162]), .I3(
        regs[130]), .S0(n46), .S1(n75), .Z(n529) );
  MUX4V2_8TH40 U366 ( .I0(regs[739]), .I1(regs[707]), .I2(regs[675]), .I3(
        regs[643]), .S0(n47), .S1(n76), .Z(n544) );
  MUX4V2_8TH40 U367 ( .I0(regs[227]), .I1(regs[195]), .I2(regs[163]), .I3(
        regs[131]), .S0(n46), .S1(n75), .Z(n539) );
  MUX4V2_8TH40 U368 ( .I0(regs[740]), .I1(regs[708]), .I2(regs[676]), .I3(
        regs[644]), .S0(n47), .S1(n76), .Z(n554) );
  MUX4V2_8TH40 U369 ( .I0(regs[228]), .I1(regs[196]), .I2(regs[164]), .I3(
        regs[132]), .S0(n47), .S1(n76), .Z(n549) );
  MUX4V2_8TH40 U370 ( .I0(regs[741]), .I1(regs[709]), .I2(regs[677]), .I3(
        regs[645]), .S0(n48), .S1(n77), .Z(n564) );
  MUX4V2_8TH40 U371 ( .I0(regs[229]), .I1(regs[197]), .I2(regs[165]), .I3(
        regs[133]), .S0(n48), .S1(n76), .Z(n559) );
  MUX4V2_8TH40 U372 ( .I0(regs[742]), .I1(regs[710]), .I2(regs[678]), .I3(
        regs[646]), .S0(n49), .S1(n77), .Z(n574) );
  MUX4V2_8TH40 U373 ( .I0(regs[230]), .I1(regs[198]), .I2(regs[166]), .I3(
        regs[134]), .S0(n48), .S1(n77), .Z(n569) );
  MUX4V2_8TH40 U374 ( .I0(regs[743]), .I1(regs[711]), .I2(regs[679]), .I3(
        regs[647]), .S0(n49), .S1(n78), .Z(n584) );
  MUX4V2_8TH40 U375 ( .I0(regs[231]), .I1(regs[199]), .I2(regs[167]), .I3(
        regs[135]), .S0(n49), .S1(n78), .Z(n579) );
  MUX4V2_8TH40 U376 ( .I0(regs[744]), .I1(regs[712]), .I2(regs[680]), .I3(
        regs[648]), .S0(n50), .S1(n79), .Z(n594) );
  MUX4V2_8TH40 U377 ( .I0(regs[232]), .I1(regs[200]), .I2(regs[168]), .I3(
        regs[136]), .S0(n50), .S1(n78), .Z(n589) );
  MUX4V2_8TH40 U378 ( .I0(regs[745]), .I1(regs[713]), .I2(regs[681]), .I3(
        regs[649]), .S0(n50), .S1(n79), .Z(n604) );
  MUX4V2_8TH40 U379 ( .I0(regs[233]), .I1(regs[201]), .I2(regs[169]), .I3(
        regs[137]), .S0(n50), .S1(n79), .Z(n599) );
  MUX4V2_8TH40 U380 ( .I0(regs[746]), .I1(regs[714]), .I2(regs[682]), .I3(
        regs[650]), .S0(n50), .S1(n80), .Z(n614) );
  MUX4V2_8TH40 U381 ( .I0(regs[234]), .I1(regs[202]), .I2(regs[170]), .I3(
        regs[138]), .S0(n51), .S1(n80), .Z(n609) );
  MUX4V2_8TH40 U382 ( .I0(regs[747]), .I1(regs[715]), .I2(regs[683]), .I3(
        regs[651]), .S0(n56), .S1(n81), .Z(n624) );
  MUX4V2_8TH40 U383 ( .I0(regs[235]), .I1(regs[203]), .I2(regs[171]), .I3(
        regs[139]), .S0(n52), .S1(n80), .Z(n619) );
  MUX4V2_8TH40 U384 ( .I0(regs[748]), .I1(regs[716]), .I2(regs[684]), .I3(
        regs[652]), .S0(n57), .S1(n81), .Z(n634) );
  MUX4V2_8TH40 U385 ( .I0(regs[236]), .I1(regs[204]), .I2(regs[172]), .I3(
        regs[140]), .S0(n58), .S1(n81), .Z(n629) );
  MUX4V2_8TH40 U386 ( .I0(regs[749]), .I1(regs[717]), .I2(regs[685]), .I3(
        regs[653]), .S0(n51), .S1(n82), .Z(n644) );
  MUX4V2_8TH40 U387 ( .I0(regs[237]), .I1(regs[205]), .I2(regs[173]), .I3(
        regs[141]), .S0(n51), .S1(n82), .Z(n639) );
  MUX4V2_8TH40 U388 ( .I0(regs[750]), .I1(regs[718]), .I2(regs[686]), .I3(
        regs[654]), .S0(n52), .S1(n82), .Z(n654) );
  MUX4V2_8TH40 U389 ( .I0(regs[238]), .I1(regs[206]), .I2(regs[174]), .I3(
        regs[142]), .S0(n51), .S1(n82), .Z(n649) );
  MUX4V2_8TH40 U390 ( .I0(regs[751]), .I1(regs[719]), .I2(regs[687]), .I3(
        regs[655]), .S0(n52), .S1(raddr1[1]), .Z(n664) );
  MUX4V2_8TH40 U391 ( .I0(regs[239]), .I1(regs[207]), .I2(regs[175]), .I3(
        regs[143]), .S0(n52), .S1(raddr1[1]), .Z(n659) );
  MUX4V2_8TH40 U392 ( .I0(regs[752]), .I1(regs[720]), .I2(regs[688]), .I3(
        regs[656]), .S0(n53), .S1(n68), .Z(n674) );
  MUX4V2_8TH40 U393 ( .I0(regs[240]), .I1(regs[208]), .I2(regs[176]), .I3(
        regs[144]), .S0(n52), .S1(n68), .Z(n669) );
  MUX4V2_8TH40 U394 ( .I0(regs[753]), .I1(regs[721]), .I2(regs[689]), .I3(
        regs[657]), .S0(n53), .S1(n69), .Z(n684) );
  MUX4V2_8TH40 U395 ( .I0(regs[241]), .I1(regs[209]), .I2(regs[177]), .I3(
        regs[145]), .S0(n53), .S1(n68), .Z(n679) );
  MUX4V2_8TH40 U396 ( .I0(regs[754]), .I1(regs[722]), .I2(regs[690]), .I3(
        regs[658]), .S0(n52), .S1(n69), .Z(n694) );
  MUX4V2_8TH40 U397 ( .I0(regs[242]), .I1(regs[210]), .I2(regs[178]), .I3(
        regs[146]), .S0(n45), .S1(n69), .Z(n689) );
  MUX4V2_8TH40 U398 ( .I0(regs[755]), .I1(regs[723]), .I2(regs[691]), .I3(
        regs[659]), .S0(n54), .S1(n70), .Z(n704) );
  MUX4V2_8TH40 U399 ( .I0(regs[243]), .I1(regs[211]), .I2(regs[179]), .I3(
        regs[147]), .S0(n46), .S1(n69), .Z(n699) );
  MUX4V2_8TH40 U400 ( .I0(regs[756]), .I1(regs[724]), .I2(regs[692]), .I3(
        regs[660]), .S0(n54), .S1(n70), .Z(n714) );
  MUX4V2_8TH40 U401 ( .I0(regs[244]), .I1(regs[212]), .I2(regs[180]), .I3(
        regs[148]), .S0(n54), .S1(n70), .Z(n709) );
  MUX4V2_8TH40 U402 ( .I0(regs[757]), .I1(regs[725]), .I2(regs[693]), .I3(
        regs[661]), .S0(n55), .S1(n71), .Z(n724) );
  MUX4V2_8TH40 U403 ( .I0(regs[245]), .I1(regs[213]), .I2(regs[181]), .I3(
        regs[149]), .S0(n56), .S1(n71), .Z(n719) );
  MUX4V2_8TH40 U404 ( .I0(regs[758]), .I1(regs[726]), .I2(regs[694]), .I3(
        regs[662]), .S0(n54), .S1(n68), .Z(n734) );
  MUX4V2_8TH40 U405 ( .I0(regs[246]), .I1(regs[214]), .I2(regs[182]), .I3(
        regs[150]), .S0(raddr1[0]), .S1(n71), .Z(n729) );
  MUX4V2_8TH40 U406 ( .I0(regs[759]), .I1(regs[727]), .I2(regs[695]), .I3(
        regs[663]), .S0(n55), .S1(n69), .Z(n744) );
  MUX4V2_8TH40 U407 ( .I0(regs[247]), .I1(regs[215]), .I2(regs[183]), .I3(
        regs[151]), .S0(n55), .S1(n74), .Z(n739) );
  MUX4V2_8TH40 U408 ( .I0(regs[760]), .I1(regs[728]), .I2(regs[696]), .I3(
        regs[664]), .S0(n56), .S1(n75), .Z(n754) );
  MUX4V2_8TH40 U409 ( .I0(regs[248]), .I1(regs[216]), .I2(regs[184]), .I3(
        regs[152]), .S0(n55), .S1(n73), .Z(n749) );
  MUX4V2_8TH40 U410 ( .I0(regs[761]), .I1(regs[729]), .I2(regs[697]), .I3(
        regs[665]), .S0(n56), .S1(n76), .Z(n764) );
  MUX4V2_8TH40 U411 ( .I0(regs[249]), .I1(regs[217]), .I2(regs[185]), .I3(
        regs[153]), .S0(n56), .S1(n77), .Z(n759) );
  MUX4V2_8TH40 U412 ( .I0(regs[762]), .I1(regs[730]), .I2(regs[698]), .I3(
        regs[666]), .S0(n57), .S1(n79), .Z(n774) );
  MUX4V2_8TH40 U413 ( .I0(regs[250]), .I1(regs[218]), .I2(regs[186]), .I3(
        regs[154]), .S0(n57), .S1(n82), .Z(n769) );
  MUX4V2_8TH40 U414 ( .I0(regs[763]), .I1(regs[731]), .I2(regs[699]), .I3(
        regs[667]), .S0(n58), .S1(n81), .Z(n784) );
  MUX4V2_8TH40 U415 ( .I0(regs[251]), .I1(regs[219]), .I2(regs[187]), .I3(
        regs[155]), .S0(n57), .S1(n80), .Z(n779) );
  MUX4V2_8TH40 U416 ( .I0(regs[764]), .I1(regs[732]), .I2(regs[700]), .I3(
        regs[668]), .S0(n58), .S1(n76), .Z(n794) );
  MUX4V2_8TH40 U417 ( .I0(regs[252]), .I1(regs[220]), .I2(regs[188]), .I3(
        regs[156]), .S0(n58), .S1(raddr1[1]), .Z(n789) );
  MUX4V2_8TH40 U418 ( .I0(regs[765]), .I1(regs[733]), .I2(regs[701]), .I3(
        regs[669]), .S0(n51), .S1(n72), .Z(n804) );
  MUX4V2_8TH40 U419 ( .I0(regs[253]), .I1(regs[221]), .I2(regs[189]), .I3(
        regs[157]), .S0(n58), .S1(n72), .Z(n799) );
  MUX4V2_8TH40 U420 ( .I0(regs[766]), .I1(regs[734]), .I2(regs[702]), .I3(
        regs[670]), .S0(n52), .S1(n73), .Z(n814) );
  MUX4V2_8TH40 U421 ( .I0(regs[254]), .I1(regs[222]), .I2(regs[190]), .I3(
        regs[158]), .S0(n45), .S1(n72), .Z(n809) );
  MUX4V2_8TH40 U422 ( .I0(regs[992]), .I1(regs[960]), .I2(regs[928]), .I3(
        regs[896]), .S0(n1), .S1(n35), .Z(n836) );
  MUX4V2_8TH40 U423 ( .I0(regs[480]), .I1(regs[448]), .I2(regs[416]), .I3(
        regs[384]), .S0(n1), .S1(n36), .Z(n831) );
  MUX4V2_8TH40 U424 ( .I0(regs[993]), .I1(regs[961]), .I2(regs[929]), .I3(
        regs[897]), .S0(n2), .S1(n31), .Z(n846) );
  MUX4V2_8TH40 U425 ( .I0(regs[481]), .I1(regs[449]), .I2(regs[417]), .I3(
        regs[385]), .S0(n1), .S1(n31), .Z(n841) );
  MUX4V2_8TH40 U426 ( .I0(regs[994]), .I1(regs[962]), .I2(regs[930]), .I3(
        regs[898]), .S0(n2), .S1(raddr2[1]), .Z(n856) );
  MUX4V2_8TH40 U427 ( .I0(regs[482]), .I1(regs[450]), .I2(regs[418]), .I3(
        regs[386]), .S0(n2), .S1(n23), .Z(n851) );
  MUX4V2_8TH40 U428 ( .I0(regs[995]), .I1(regs[963]), .I2(regs[931]), .I3(
        regs[899]), .S0(n3), .S1(n31), .Z(n866) );
  MUX4V2_8TH40 U429 ( .I0(regs[483]), .I1(regs[451]), .I2(regs[419]), .I3(
        regs[387]), .S0(n3), .S1(n24), .Z(n861) );
  MUX4V2_8TH40 U430 ( .I0(regs[996]), .I1(regs[964]), .I2(regs[932]), .I3(
        regs[900]), .S0(n4), .S1(n31), .Z(n876) );
  MUX4V2_8TH40 U431 ( .I0(regs[484]), .I1(regs[452]), .I2(regs[420]), .I3(
        regs[388]), .S0(n3), .S1(n31), .Z(n871) );
  MUX4V2_8TH40 U432 ( .I0(regs[997]), .I1(regs[965]), .I2(regs[933]), .I3(
        regs[901]), .S0(n4), .S1(n32), .Z(n886) );
  MUX4V2_8TH40 U433 ( .I0(regs[485]), .I1(regs[453]), .I2(regs[421]), .I3(
        regs[389]), .S0(n4), .S1(n32), .Z(n881) );
  MUX4V2_8TH40 U434 ( .I0(regs[998]), .I1(regs[966]), .I2(regs[934]), .I3(
        regs[902]), .S0(n5), .S1(n33), .Z(n896) );
  MUX4V2_8TH40 U435 ( .I0(regs[486]), .I1(regs[454]), .I2(regs[422]), .I3(
        regs[390]), .S0(n4), .S1(n32), .Z(n891) );
  MUX4V2_8TH40 U436 ( .I0(regs[999]), .I1(regs[967]), .I2(regs[935]), .I3(
        regs[903]), .S0(n5), .S1(n33), .Z(n906) );
  MUX4V2_8TH40 U437 ( .I0(regs[487]), .I1(regs[455]), .I2(regs[423]), .I3(
        regs[391]), .S0(n5), .S1(n33), .Z(n901) );
  MUX4V2_8TH40 U438 ( .I0(regs[1000]), .I1(regs[968]), .I2(regs[936]), .I3(
        regs[904]), .S0(n6), .S1(n34), .Z(n916) );
  MUX4V2_8TH40 U439 ( .I0(regs[488]), .I1(regs[456]), .I2(regs[424]), .I3(
        regs[392]), .S0(n6), .S1(n34), .Z(n911) );
  MUX4V2_8TH40 U440 ( .I0(regs[1001]), .I1(regs[969]), .I2(regs[937]), .I3(
        regs[905]), .S0(n7), .S1(n35), .Z(n926) );
  MUX4V2_8TH40 U441 ( .I0(regs[489]), .I1(regs[457]), .I2(regs[425]), .I3(
        regs[393]), .S0(n6), .S1(n34), .Z(n921) );
  MUX4V2_8TH40 U442 ( .I0(regs[1002]), .I1(regs[970]), .I2(regs[938]), .I3(
        regs[906]), .S0(n7), .S1(n35), .Z(n936) );
  MUX4V2_8TH40 U443 ( .I0(regs[490]), .I1(regs[458]), .I2(regs[426]), .I3(
        regs[394]), .S0(n7), .S1(n35), .Z(n931) );
  MUX4V2_8TH40 U444 ( .I0(regs[1003]), .I1(regs[971]), .I2(regs[939]), .I3(
        regs[907]), .S0(n8), .S1(n36), .Z(n946) );
  MUX4V2_8TH40 U445 ( .I0(regs[491]), .I1(regs[459]), .I2(regs[427]), .I3(
        regs[395]), .S0(n8), .S1(n35), .Z(n941) );
  MUX4V2_8TH40 U446 ( .I0(regs[1004]), .I1(regs[972]), .I2(regs[940]), .I3(
        regs[908]), .S0(n8), .S1(n36), .Z(n956) );
  MUX4V2_8TH40 U447 ( .I0(regs[492]), .I1(regs[460]), .I2(regs[428]), .I3(
        regs[396]), .S0(n8), .S1(n36), .Z(n951) );
  MUX4V2_8TH40 U448 ( .I0(regs[1005]), .I1(regs[973]), .I2(regs[941]), .I3(
        regs[909]), .S0(n9), .S1(n31), .Z(n966) );
  MUX4V2_8TH40 U449 ( .I0(regs[493]), .I1(regs[461]), .I2(regs[429]), .I3(
        regs[397]), .S0(n9), .S1(n32), .Z(n961) );
  MUX4V2_8TH40 U450 ( .I0(regs[1006]), .I1(regs[974]), .I2(regs[942]), .I3(
        regs[910]), .S0(n10), .S1(raddr2[1]), .Z(n976) );
  MUX4V2_8TH40 U451 ( .I0(regs[494]), .I1(regs[462]), .I2(regs[430]), .I3(
        regs[398]), .S0(n9), .S1(n25), .Z(n971) );
  MUX4V2_8TH40 U452 ( .I0(regs[1007]), .I1(regs[975]), .I2(regs[943]), .I3(
        regs[911]), .S0(n10), .S1(raddr2[1]), .Z(n986) );
  MUX4V2_8TH40 U453 ( .I0(regs[495]), .I1(regs[463]), .I2(regs[431]), .I3(
        regs[399]), .S0(n10), .S1(raddr2[1]), .Z(n981) );
  MUX4V2_8TH40 U454 ( .I0(regs[1008]), .I1(regs[976]), .I2(regs[944]), .I3(
        regs[912]), .S0(n11), .S1(n23), .Z(n996) );
  MUX4V2_8TH40 U455 ( .I0(regs[496]), .I1(regs[464]), .I2(regs[432]), .I3(
        regs[400]), .S0(n11), .S1(n23), .Z(n991) );
  MUX4V2_8TH40 U456 ( .I0(regs[1009]), .I1(regs[977]), .I2(regs[945]), .I3(
        regs[913]), .S0(n12), .S1(n24), .Z(n1006) );
  MUX4V2_8TH40 U457 ( .I0(regs[497]), .I1(regs[465]), .I2(regs[433]), .I3(
        regs[401]), .S0(n11), .S1(n23), .Z(n1001) );
  MUX4V2_8TH40 U458 ( .I0(regs[1010]), .I1(regs[978]), .I2(regs[946]), .I3(
        regs[914]), .S0(n12), .S1(n24), .Z(n1016) );
  MUX4V2_8TH40 U459 ( .I0(regs[498]), .I1(regs[466]), .I2(regs[434]), .I3(
        regs[402]), .S0(n12), .S1(n24), .Z(n1011) );
  MUX4V2_8TH40 U460 ( .I0(regs[1011]), .I1(regs[979]), .I2(regs[947]), .I3(
        regs[915]), .S0(n12), .S1(n25), .Z(n1026) );
  MUX4V2_8TH40 U461 ( .I0(regs[499]), .I1(regs[467]), .I2(regs[435]), .I3(
        regs[403]), .S0(n12), .S1(n25), .Z(n1021) );
  MUX4V2_8TH40 U462 ( .I0(regs[1012]), .I1(regs[980]), .I2(regs[948]), .I3(
        regs[916]), .S0(n13), .S1(n26), .Z(n1036) );
  MUX4V2_8TH40 U463 ( .I0(regs[500]), .I1(regs[468]), .I2(regs[436]), .I3(
        regs[404]), .S0(n14), .S1(n25), .Z(n1031) );
  MUX4V2_8TH40 U464 ( .I0(regs[1013]), .I1(regs[981]), .I2(regs[949]), .I3(
        regs[917]), .S0(n2), .S1(n26), .Z(n1046) );
  MUX4V2_8TH40 U465 ( .I0(regs[501]), .I1(regs[469]), .I2(regs[437]), .I3(
        regs[405]), .S0(n4), .S1(n26), .Z(n1041) );
  MUX4V2_8TH40 U466 ( .I0(regs[1014]), .I1(regs[982]), .I2(regs[950]), .I3(
        regs[918]), .S0(n8), .S1(n27), .Z(n1056) );
  MUX4V2_8TH40 U467 ( .I0(regs[502]), .I1(regs[470]), .I2(regs[438]), .I3(
        regs[406]), .S0(n3), .S1(n26), .Z(n1051) );
  MUX4V2_8TH40 U468 ( .I0(regs[1015]), .I1(regs[983]), .I2(regs[951]), .I3(
        regs[919]), .S0(n11), .S1(n27), .Z(n1066) );
  MUX4V2_8TH40 U469 ( .I0(regs[503]), .I1(regs[471]), .I2(regs[439]), .I3(
        regs[407]), .S0(n12), .S1(n27), .Z(n1061) );
  MUX4V2_8TH40 U470 ( .I0(regs[1016]), .I1(regs[984]), .I2(regs[952]), .I3(
        regs[920]), .S0(n8), .S1(n28), .Z(n1076) );
  MUX4V2_8TH40 U471 ( .I0(regs[504]), .I1(regs[472]), .I2(regs[440]), .I3(
        regs[408]), .S0(n11), .S1(n28), .Z(n1071) );
  MUX4V2_8TH40 U472 ( .I0(regs[1017]), .I1(regs[985]), .I2(regs[953]), .I3(
        regs[921]), .S0(n12), .S1(n29), .Z(n1086) );
  MUX4V2_8TH40 U473 ( .I0(regs[505]), .I1(regs[473]), .I2(regs[441]), .I3(
        regs[409]), .S0(n13), .S1(n28), .Z(n1081) );
  MUX4V2_8TH40 U474 ( .I0(regs[1018]), .I1(regs[986]), .I2(regs[954]), .I3(
        regs[922]), .S0(n13), .S1(n29), .Z(n1096) );
  MUX4V2_8TH40 U475 ( .I0(regs[506]), .I1(regs[474]), .I2(regs[442]), .I3(
        regs[410]), .S0(n13), .S1(n29), .Z(n1091) );
  MUX4V2_8TH40 U476 ( .I0(regs[1019]), .I1(regs[987]), .I2(regs[955]), .I3(
        regs[923]), .S0(n14), .S1(n30), .Z(n1106) );
  MUX4V2_8TH40 U477 ( .I0(regs[507]), .I1(regs[475]), .I2(regs[443]), .I3(
        regs[411]), .S0(n13), .S1(n30), .Z(n1101) );
  MUX4V2_8TH40 U478 ( .I0(regs[1020]), .I1(regs[988]), .I2(regs[956]), .I3(
        regs[924]), .S0(n14), .S1(n30), .Z(n1116) );
  MUX4V2_8TH40 U479 ( .I0(regs[508]), .I1(regs[476]), .I2(regs[444]), .I3(
        regs[412]), .S0(n14), .S1(n30), .Z(n1111) );
  MUX4V2_8TH40 U480 ( .I0(regs[1021]), .I1(regs[989]), .I2(regs[957]), .I3(
        regs[925]), .S0(raddr2[0]), .S1(n30), .Z(n1126) );
  MUX4V2_8TH40 U481 ( .I0(regs[509]), .I1(regs[477]), .I2(regs[445]), .I3(
        regs[413]), .S0(raddr2[0]), .S1(n33), .Z(n1121) );
  MUX4V2_8TH40 U482 ( .I0(regs[510]), .I1(regs[478]), .I2(regs[446]), .I3(
        regs[414]), .S0(raddr2[0]), .S1(n34), .Z(n1131) );
  MUX4V2_8TH40 U483 ( .I0(regs[992]), .I1(regs[960]), .I2(regs[928]), .I3(
        regs[896]), .S0(n45), .S1(n74), .Z(n100) );
  MUX4V2_8TH40 U484 ( .I0(regs[480]), .I1(regs[448]), .I2(regs[416]), .I3(
        regs[384]), .S0(n45), .S1(n74), .Z(n95) );
  MUX4V2_8TH40 U485 ( .I0(regs[993]), .I1(regs[961]), .I2(regs[929]), .I3(
        regs[897]), .S0(n46), .S1(n74), .Z(n110) );
  MUX4V2_8TH40 U486 ( .I0(regs[481]), .I1(regs[449]), .I2(regs[417]), .I3(
        regs[385]), .S0(n45), .S1(n74), .Z(n105) );
  MUX4V2_8TH40 U487 ( .I0(regs[994]), .I1(regs[962]), .I2(regs[930]), .I3(
        regs[898]), .S0(n46), .S1(n75), .Z(n536) );
  MUX4V2_8TH40 U488 ( .I0(regs[482]), .I1(regs[450]), .I2(regs[418]), .I3(
        regs[386]), .S0(n46), .S1(n75), .Z(n531) );
  MUX4V2_8TH40 U489 ( .I0(regs[995]), .I1(regs[963]), .I2(regs[931]), .I3(
        regs[899]), .S0(n47), .S1(n76), .Z(n546) );
  MUX4V2_8TH40 U490 ( .I0(regs[483]), .I1(regs[451]), .I2(regs[419]), .I3(
        regs[387]), .S0(n47), .S1(n75), .Z(n541) );
  MUX4V2_8TH40 U491 ( .I0(regs[996]), .I1(regs[964]), .I2(regs[932]), .I3(
        regs[900]), .S0(n48), .S1(n76), .Z(n556) );
  MUX4V2_8TH40 U492 ( .I0(regs[484]), .I1(regs[452]), .I2(regs[420]), .I3(
        regs[388]), .S0(n47), .S1(n76), .Z(n551) );
  MUX4V2_8TH40 U493 ( .I0(regs[997]), .I1(regs[965]), .I2(regs[933]), .I3(
        regs[901]), .S0(n48), .S1(n77), .Z(n566) );
  MUX4V2_8TH40 U494 ( .I0(regs[485]), .I1(regs[453]), .I2(regs[421]), .I3(
        regs[389]), .S0(n48), .S1(n77), .Z(n561) );
  MUX4V2_8TH40 U495 ( .I0(regs[998]), .I1(regs[966]), .I2(regs[934]), .I3(
        regs[902]), .S0(n49), .S1(n78), .Z(n576) );
  MUX4V2_8TH40 U496 ( .I0(regs[486]), .I1(regs[454]), .I2(regs[422]), .I3(
        regs[390]), .S0(n48), .S1(n77), .Z(n571) );
  MUX4V2_8TH40 U497 ( .I0(regs[999]), .I1(regs[967]), .I2(regs[935]), .I3(
        regs[903]), .S0(n49), .S1(n78), .Z(n586) );
  MUX4V2_8TH40 U498 ( .I0(regs[487]), .I1(regs[455]), .I2(regs[423]), .I3(
        regs[391]), .S0(n49), .S1(n78), .Z(n581) );
  MUX4V2_8TH40 U499 ( .I0(regs[1000]), .I1(regs[968]), .I2(regs[936]), .I3(
        regs[904]), .S0(n50), .S1(n79), .Z(n596) );
  MUX4V2_8TH40 U500 ( .I0(regs[488]), .I1(regs[456]), .I2(regs[424]), .I3(
        regs[392]), .S0(n50), .S1(n79), .Z(n591) );
  MUX4V2_8TH40 U501 ( .I0(regs[1001]), .I1(regs[969]), .I2(regs[937]), .I3(
        regs[905]), .S0(n45), .S1(n80), .Z(n606) );
  MUX4V2_8TH40 U502 ( .I0(regs[489]), .I1(regs[457]), .I2(regs[425]), .I3(
        regs[393]), .S0(n50), .S1(n79), .Z(n601) );
  MUX4V2_8TH40 U503 ( .I0(regs[1002]), .I1(regs[970]), .I2(regs[938]), .I3(
        regs[906]), .S0(n46), .S1(n80), .Z(n616) );
  MUX4V2_8TH40 U504 ( .I0(regs[490]), .I1(regs[458]), .I2(regs[426]), .I3(
        regs[394]), .S0(n47), .S1(n80), .Z(n611) );
  MUX4V2_8TH40 U505 ( .I0(regs[1003]), .I1(regs[971]), .I2(regs[939]), .I3(
        regs[907]), .S0(n46), .S1(n81), .Z(n626) );
  MUX4V2_8TH40 U506 ( .I0(regs[491]), .I1(regs[459]), .I2(regs[427]), .I3(
        regs[395]), .S0(n47), .S1(n80), .Z(n621) );
  MUX4V2_8TH40 U507 ( .I0(regs[1004]), .I1(regs[972]), .I2(regs[940]), .I3(
        regs[908]), .S0(n48), .S1(n81), .Z(n636) );
  MUX4V2_8TH40 U508 ( .I0(regs[492]), .I1(regs[460]), .I2(regs[428]), .I3(
        regs[396]), .S0(n53), .S1(n81), .Z(n631) );
  MUX4V2_8TH40 U509 ( .I0(regs[1005]), .I1(regs[973]), .I2(regs[941]), .I3(
        regs[909]), .S0(n51), .S1(n82), .Z(n646) );
  MUX4V2_8TH40 U510 ( .I0(regs[493]), .I1(regs[461]), .I2(regs[429]), .I3(
        regs[397]), .S0(n51), .S1(n82), .Z(n641) );
  MUX4V2_8TH40 U511 ( .I0(regs[1006]), .I1(regs[974]), .I2(regs[942]), .I3(
        regs[910]), .S0(n52), .S1(raddr1[1]), .Z(n656) );
  MUX4V2_8TH40 U512 ( .I0(regs[494]), .I1(regs[462]), .I2(regs[430]), .I3(
        regs[398]), .S0(n51), .S1(n82), .Z(n651) );
  MUX4V2_8TH40 U513 ( .I0(regs[1007]), .I1(regs[975]), .I2(regs[943]), .I3(
        regs[911]), .S0(n52), .S1(raddr1[1]), .Z(n666) );
  MUX4V2_8TH40 U514 ( .I0(regs[495]), .I1(regs[463]), .I2(regs[431]), .I3(
        regs[399]), .S0(n52), .S1(raddr1[1]), .Z(n661) );
  MUX4V2_8TH40 U515 ( .I0(regs[496]), .I1(regs[464]), .I2(regs[432]), .I3(
        regs[400]), .S0(n53), .S1(n68), .Z(n671) );
  MUX4V2_8TH40 U516 ( .I0(regs[497]), .I1(regs[465]), .I2(regs[433]), .I3(
        regs[401]), .S0(n53), .S1(n68), .Z(n681) );
  MUX4V2_8TH40 U517 ( .I0(regs[498]), .I1(regs[466]), .I2(regs[434]), .I3(
        regs[402]), .S0(n47), .S1(n69), .Z(n691) );
  MUX4V2_8TH40 U518 ( .I0(regs[499]), .I1(regs[467]), .I2(regs[435]), .I3(
        regs[403]), .S0(n48), .S1(n70), .Z(n701) );
  MUX4V2_8TH40 U519 ( .I0(regs[500]), .I1(regs[468]), .I2(regs[436]), .I3(
        regs[404]), .S0(n54), .S1(n70), .Z(n711) );
  MUX4V2_8TH40 U520 ( .I0(regs[501]), .I1(regs[469]), .I2(regs[437]), .I3(
        regs[405]), .S0(n49), .S1(n71), .Z(n721) );
  MUX4V2_8TH40 U521 ( .I0(regs[502]), .I1(regs[470]), .I2(regs[438]), .I3(
        regs[406]), .S0(n50), .S1(n71), .Z(n731) );
  MUX4V2_8TH40 U522 ( .I0(regs[503]), .I1(regs[471]), .I2(regs[439]), .I3(
        regs[407]), .S0(n55), .S1(n75), .Z(n741) );
  MUX4V2_8TH40 U523 ( .I0(regs[504]), .I1(regs[472]), .I2(regs[440]), .I3(
        regs[408]), .S0(n56), .S1(n70), .Z(n751) );
  MUX4V2_8TH40 U524 ( .I0(regs[505]), .I1(regs[473]), .I2(regs[441]), .I3(
        regs[409]), .S0(n56), .S1(n71), .Z(n761) );
  MUX4V2_8TH40 U525 ( .I0(regs[506]), .I1(regs[474]), .I2(regs[442]), .I3(
        regs[410]), .S0(n57), .S1(n81), .Z(n771) );
  MUX4V2_8TH40 U526 ( .I0(regs[507]), .I1(regs[475]), .I2(regs[443]), .I3(
        regs[411]), .S0(n57), .S1(n68), .Z(n781) );
  MUX4V2_8TH40 U527 ( .I0(regs[508]), .I1(regs[476]), .I2(regs[444]), .I3(
        regs[412]), .S0(n58), .S1(n69), .Z(n791) );
  MUX4V2_8TH40 U528 ( .I0(regs[509]), .I1(regs[477]), .I2(regs[445]), .I3(
        regs[413]), .S0(n46), .S1(n72), .Z(n801) );
  MUX4V2_8TH40 U529 ( .I0(regs[510]), .I1(regs[478]), .I2(regs[446]), .I3(
        regs[414]), .S0(n57), .S1(n72), .Z(n811) );
  MUX4V2_8TH40 U530 ( .I0(regs[767]), .I1(regs[735]), .I2(regs[703]), .I3(
        regs[671]), .S0(n6), .S1(n29), .Z(n1144) );
  MUX4V2_8TH40 U531 ( .I0(regs[255]), .I1(regs[223]), .I2(regs[191]), .I3(
        regs[159]), .S0(n9), .S1(n30), .Z(n1139) );
  MUX4V2_8TH40 U532 ( .I0(regs[767]), .I1(regs[735]), .I2(regs[703]), .I3(
        regs[671]), .S0(raddr1[0]), .S1(n73), .Z(n824) );
  MUX4V2_8TH40 U533 ( .I0(regs[255]), .I1(regs[223]), .I2(regs[191]), .I3(
        regs[159]), .S0(raddr1[0]), .S1(n73), .Z(n819) );
  MUX4V2_8TH40 U534 ( .I0(regs[1022]), .I1(regs[990]), .I2(regs[958]), .I3(
        regs[926]), .S0(n10), .S1(n33), .Z(n1136) );
  MUX4V2_8TH40 U535 ( .I0(regs[1023]), .I1(regs[991]), .I2(regs[959]), .I3(
        regs[927]), .S0(n1), .S1(n34), .Z(n1146) );
  MUX4V2_8TH40 U536 ( .I0(regs[511]), .I1(regs[479]), .I2(regs[447]), .I3(
        regs[415]), .S0(n2), .S1(n35), .Z(n1141) );
  MUX4V2_8TH40 U537 ( .I0(regs[511]), .I1(regs[479]), .I2(regs[447]), .I3(
        regs[415]), .S0(raddr1[0]), .S1(n73), .Z(n821) );
  MUX4V2_8TH40 U538 ( .I0(regs[864]), .I1(regs[832]), .I2(regs[800]), .I3(
        regs[768]), .S0(n1), .S1(raddr2[1]), .Z(n835) );
  MUX4V2_8TH40 U539 ( .I0(regs[352]), .I1(regs[320]), .I2(regs[288]), .I3(
        regs[256]), .S0(n1), .S1(n36), .Z(n830) );
  MUX4V2_8TH40 U540 ( .I0(regs[865]), .I1(regs[833]), .I2(regs[801]), .I3(
        regs[769]), .S0(n2), .S1(n23), .Z(n845) );
  MUX4V2_8TH40 U541 ( .I0(regs[353]), .I1(regs[321]), .I2(regs[289]), .I3(
        regs[257]), .S0(n1), .S1(n24), .Z(n840) );
  MUX4V2_8TH40 U542 ( .I0(regs[866]), .I1(regs[834]), .I2(regs[802]), .I3(
        regs[770]), .S0(n2), .S1(n27), .Z(n855) );
  MUX4V2_8TH40 U543 ( .I0(regs[354]), .I1(regs[322]), .I2(regs[290]), .I3(
        regs[258]), .S0(n2), .S1(n28), .Z(n850) );
  MUX4V2_8TH40 U544 ( .I0(regs[867]), .I1(regs[835]), .I2(regs[803]), .I3(
        regs[771]), .S0(n3), .S1(n31), .Z(n865) );
  MUX4V2_8TH40 U545 ( .I0(regs[355]), .I1(regs[323]), .I2(regs[291]), .I3(
        regs[259]), .S0(n3), .S1(n31), .Z(n860) );
  MUX4V2_8TH40 U546 ( .I0(regs[868]), .I1(regs[836]), .I2(regs[804]), .I3(
        regs[772]), .S0(n3), .S1(n31), .Z(n875) );
  MUX4V2_8TH40 U547 ( .I0(regs[356]), .I1(regs[324]), .I2(regs[292]), .I3(
        regs[260]), .S0(n3), .S1(n31), .Z(n870) );
  MUX4V2_8TH40 U548 ( .I0(regs[869]), .I1(regs[837]), .I2(regs[805]), .I3(
        regs[773]), .S0(n4), .S1(n32), .Z(n885) );
  MUX4V2_8TH40 U549 ( .I0(regs[357]), .I1(regs[325]), .I2(regs[293]), .I3(
        regs[261]), .S0(n4), .S1(n32), .Z(n880) );
  MUX4V2_8TH40 U550 ( .I0(regs[870]), .I1(regs[838]), .I2(regs[806]), .I3(
        regs[774]), .S0(n5), .S1(n32), .Z(n895) );
  MUX4V2_8TH40 U551 ( .I0(regs[358]), .I1(regs[326]), .I2(regs[294]), .I3(
        regs[262]), .S0(n4), .S1(n32), .Z(n890) );
  MUX4V2_8TH40 U552 ( .I0(regs[871]), .I1(regs[839]), .I2(regs[807]), .I3(
        regs[775]), .S0(n5), .S1(n33), .Z(n905) );
  MUX4V2_8TH40 U553 ( .I0(regs[359]), .I1(regs[327]), .I2(regs[295]), .I3(
        regs[263]), .S0(n5), .S1(n33), .Z(n900) );
  MUX4V2_8TH40 U554 ( .I0(regs[872]), .I1(regs[840]), .I2(regs[808]), .I3(
        regs[776]), .S0(n6), .S1(n34), .Z(n915) );
  MUX4V2_8TH40 U555 ( .I0(regs[360]), .I1(regs[328]), .I2(regs[296]), .I3(
        regs[264]), .S0(n6), .S1(n33), .Z(n910) );
  MUX4V2_8TH40 U556 ( .I0(regs[873]), .I1(regs[841]), .I2(regs[809]), .I3(
        regs[777]), .S0(n7), .S1(n34), .Z(n925) );
  MUX4V2_8TH40 U557 ( .I0(regs[361]), .I1(regs[329]), .I2(regs[297]), .I3(
        regs[265]), .S0(n6), .S1(n34), .Z(n920) );
  MUX4V2_8TH40 U558 ( .I0(regs[874]), .I1(regs[842]), .I2(regs[810]), .I3(
        regs[778]), .S0(n7), .S1(n35), .Z(n935) );
  MUX4V2_8TH40 U559 ( .I0(regs[362]), .I1(regs[330]), .I2(regs[298]), .I3(
        regs[266]), .S0(n7), .S1(n35), .Z(n930) );
  MUX4V2_8TH40 U560 ( .I0(regs[875]), .I1(regs[843]), .I2(regs[811]), .I3(
        regs[779]), .S0(n8), .S1(n36), .Z(n945) );
  MUX4V2_8TH40 U561 ( .I0(regs[363]), .I1(regs[331]), .I2(regs[299]), .I3(
        regs[267]), .S0(n7), .S1(n35), .Z(n940) );
  MUX4V2_8TH40 U562 ( .I0(regs[876]), .I1(regs[844]), .I2(regs[812]), .I3(
        regs[780]), .S0(n8), .S1(n36), .Z(n955) );
  MUX4V2_8TH40 U563 ( .I0(regs[364]), .I1(regs[332]), .I2(regs[300]), .I3(
        regs[268]), .S0(n8), .S1(n36), .Z(n950) );
  MUX4V2_8TH40 U564 ( .I0(regs[877]), .I1(regs[845]), .I2(regs[813]), .I3(
        regs[781]), .S0(n9), .S1(n26), .Z(n965) );
  MUX4V2_8TH40 U565 ( .I0(regs[365]), .I1(regs[333]), .I2(regs[301]), .I3(
        regs[269]), .S0(n9), .S1(n36), .Z(n960) );
  MUX4V2_8TH40 U566 ( .I0(regs[878]), .I1(regs[846]), .I2(regs[814]), .I3(
        regs[782]), .S0(n10), .S1(n29), .Z(n975) );
  MUX4V2_8TH40 U567 ( .I0(regs[366]), .I1(regs[334]), .I2(regs[302]), .I3(
        regs[270]), .S0(n9), .S1(n30), .Z(n970) );
  MUX4V2_8TH40 U568 ( .I0(regs[879]), .I1(regs[847]), .I2(regs[815]), .I3(
        regs[783]), .S0(n10), .S1(raddr2[1]), .Z(n985) );
  MUX4V2_8TH40 U569 ( .I0(regs[367]), .I1(regs[335]), .I2(regs[303]), .I3(
        regs[271]), .S0(n10), .S1(raddr2[1]), .Z(n980) );
  MUX4V2_8TH40 U570 ( .I0(regs[880]), .I1(regs[848]), .I2(regs[816]), .I3(
        regs[784]), .S0(n11), .S1(n23), .Z(n995) );
  MUX4V2_8TH40 U571 ( .I0(regs[368]), .I1(regs[336]), .I2(regs[304]), .I3(
        regs[272]), .S0(n11), .S1(n23), .Z(n990) );
  MUX4V2_8TH40 U572 ( .I0(regs[881]), .I1(regs[849]), .I2(regs[817]), .I3(
        regs[785]), .S0(n11), .S1(n24), .Z(n1005) );
  MUX4V2_8TH40 U573 ( .I0(regs[369]), .I1(regs[337]), .I2(regs[305]), .I3(
        regs[273]), .S0(n11), .S1(n23), .Z(n1000) );
  MUX4V2_8TH40 U574 ( .I0(regs[882]), .I1(regs[850]), .I2(regs[818]), .I3(
        regs[786]), .S0(n12), .S1(n24), .Z(n1015) );
  MUX4V2_8TH40 U575 ( .I0(regs[370]), .I1(regs[338]), .I2(regs[306]), .I3(
        regs[274]), .S0(n12), .S1(n24), .Z(n1010) );
  MUX4V2_8TH40 U576 ( .I0(regs[883]), .I1(regs[851]), .I2(regs[819]), .I3(
        regs[787]), .S0(n9), .S1(n25), .Z(n1025) );
  MUX4V2_8TH40 U577 ( .I0(regs[371]), .I1(regs[339]), .I2(regs[307]), .I3(
        regs[275]), .S0(n12), .S1(n25), .Z(n1020) );
  MUX4V2_8TH40 U578 ( .I0(regs[884]), .I1(regs[852]), .I2(regs[820]), .I3(
        regs[788]), .S0(n9), .S1(n25), .Z(n1035) );
  MUX4V2_8TH40 U579 ( .I0(regs[372]), .I1(regs[340]), .I2(regs[308]), .I3(
        regs[276]), .S0(n4), .S1(n25), .Z(n1030) );
  MUX4V2_8TH40 U580 ( .I0(regs[885]), .I1(regs[853]), .I2(regs[821]), .I3(
        regs[789]), .S0(raddr2[0]), .S1(n26), .Z(n1045) );
  MUX4V2_8TH40 U581 ( .I0(regs[373]), .I1(regs[341]), .I2(regs[309]), .I3(
        regs[277]), .S0(n5), .S1(n26), .Z(n1040) );
  MUX4V2_8TH40 U582 ( .I0(regs[886]), .I1(regs[854]), .I2(regs[822]), .I3(
        regs[790]), .S0(n13), .S1(n27), .Z(n1055) );
  MUX4V2_8TH40 U583 ( .I0(regs[374]), .I1(regs[342]), .I2(regs[310]), .I3(
        regs[278]), .S0(n6), .S1(n26), .Z(n1050) );
  MUX4V2_8TH40 U584 ( .I0(regs[887]), .I1(regs[855]), .I2(regs[823]), .I3(
        regs[791]), .S0(n14), .S1(n27), .Z(n1065) );
  MUX4V2_8TH40 U585 ( .I0(regs[375]), .I1(regs[343]), .I2(regs[311]), .I3(
        regs[279]), .S0(n4), .S1(n27), .Z(n1060) );
  MUX4V2_8TH40 U586 ( .I0(regs[888]), .I1(regs[856]), .I2(regs[824]), .I3(
        regs[792]), .S0(n14), .S1(n28), .Z(n1075) );
  MUX4V2_8TH40 U587 ( .I0(regs[376]), .I1(regs[344]), .I2(regs[312]), .I3(
        regs[280]), .S0(n3), .S1(n28), .Z(n1070) );
  MUX4V2_8TH40 U588 ( .I0(regs[889]), .I1(regs[857]), .I2(regs[825]), .I3(
        regs[793]), .S0(n6), .S1(n29), .Z(n1085) );
  MUX4V2_8TH40 U589 ( .I0(regs[377]), .I1(regs[345]), .I2(regs[313]), .I3(
        regs[281]), .S0(n4), .S1(n28), .Z(n1080) );
  MUX4V2_8TH40 U590 ( .I0(regs[890]), .I1(regs[858]), .I2(regs[826]), .I3(
        regs[794]), .S0(n13), .S1(n29), .Z(n1095) );
  MUX4V2_8TH40 U591 ( .I0(regs[378]), .I1(regs[346]), .I2(regs[314]), .I3(
        regs[282]), .S0(n13), .S1(n29), .Z(n1090) );
  MUX4V2_8TH40 U592 ( .I0(regs[891]), .I1(regs[859]), .I2(regs[827]), .I3(
        regs[795]), .S0(n14), .S1(n30), .Z(n1105) );
  MUX4V2_8TH40 U593 ( .I0(regs[379]), .I1(regs[347]), .I2(regs[315]), .I3(
        regs[283]), .S0(n13), .S1(n29), .Z(n1100) );
  MUX4V2_8TH40 U594 ( .I0(regs[892]), .I1(regs[860]), .I2(regs[828]), .I3(
        regs[796]), .S0(n14), .S1(n30), .Z(n1115) );
  MUX4V2_8TH40 U595 ( .I0(regs[380]), .I1(regs[348]), .I2(regs[316]), .I3(
        regs[284]), .S0(n14), .S1(n30), .Z(n1110) );
  MUX4V2_8TH40 U596 ( .I0(regs[893]), .I1(regs[861]), .I2(regs[829]), .I3(
        regs[797]), .S0(raddr2[0]), .S1(n35), .Z(n1125) );
  MUX4V2_8TH40 U597 ( .I0(regs[381]), .I1(regs[349]), .I2(regs[317]), .I3(
        regs[285]), .S0(raddr2[0]), .S1(n36), .Z(n1120) );
  MUX4V2_8TH40 U598 ( .I0(regs[894]), .I1(regs[862]), .I2(regs[830]), .I3(
        regs[798]), .S0(raddr2[0]), .S1(n28), .Z(n1135) );
  MUX4V2_8TH40 U599 ( .I0(regs[382]), .I1(regs[350]), .I2(regs[318]), .I3(
        regs[286]), .S0(raddr2[0]), .S1(raddr2[1]), .Z(n1130) );
  MUX4V2_8TH40 U600 ( .I0(regs[864]), .I1(regs[832]), .I2(regs[800]), .I3(
        regs[768]), .S0(n45), .S1(n74), .Z(n99) );
  MUX4V2_8TH40 U601 ( .I0(regs[352]), .I1(regs[320]), .I2(regs[288]), .I3(
        regs[256]), .S0(n45), .S1(n73), .Z(n94) );
  MUX4V2_8TH40 U602 ( .I0(regs[865]), .I1(regs[833]), .I2(regs[801]), .I3(
        regs[769]), .S0(n46), .S1(n74), .Z(n109) );
  MUX4V2_8TH40 U603 ( .I0(regs[353]), .I1(regs[321]), .I2(regs[289]), .I3(
        regs[257]), .S0(n45), .S1(n74), .Z(n104) );
  MUX4V2_8TH40 U604 ( .I0(regs[866]), .I1(regs[834]), .I2(regs[802]), .I3(
        regs[770]), .S0(n46), .S1(n75), .Z(n535) );
  MUX4V2_8TH40 U605 ( .I0(regs[354]), .I1(regs[322]), .I2(regs[290]), .I3(
        regs[258]), .S0(n46), .S1(n75), .Z(n530) );
  MUX4V2_8TH40 U606 ( .I0(regs[867]), .I1(regs[835]), .I2(regs[803]), .I3(
        regs[771]), .S0(n47), .S1(n76), .Z(n545) );
  MUX4V2_8TH40 U607 ( .I0(regs[355]), .I1(regs[323]), .I2(regs[291]), .I3(
        regs[259]), .S0(n47), .S1(n75), .Z(n540) );
  MUX4V2_8TH40 U608 ( .I0(regs[868]), .I1(regs[836]), .I2(regs[804]), .I3(
        regs[772]), .S0(n47), .S1(n76), .Z(n555) );
  MUX4V2_8TH40 U609 ( .I0(regs[356]), .I1(regs[324]), .I2(regs[292]), .I3(
        regs[260]), .S0(n47), .S1(n76), .Z(n550) );
  MUX4V2_8TH40 U610 ( .I0(regs[869]), .I1(regs[837]), .I2(regs[805]), .I3(
        regs[773]), .S0(n48), .S1(n77), .Z(n565) );
  MUX4V2_8TH40 U611 ( .I0(regs[357]), .I1(regs[325]), .I2(regs[293]), .I3(
        regs[261]), .S0(n48), .S1(n77), .Z(n560) );
  MUX4V2_8TH40 U612 ( .I0(regs[870]), .I1(regs[838]), .I2(regs[806]), .I3(
        regs[774]), .S0(n49), .S1(n77), .Z(n575) );
  MUX4V2_8TH40 U613 ( .I0(regs[358]), .I1(regs[326]), .I2(regs[294]), .I3(
        regs[262]), .S0(n48), .S1(n77), .Z(n570) );
  MUX4V2_8TH40 U614 ( .I0(regs[871]), .I1(regs[839]), .I2(regs[807]), .I3(
        regs[775]), .S0(n49), .S1(n78), .Z(n585) );
  MUX4V2_8TH40 U615 ( .I0(regs[359]), .I1(regs[327]), .I2(regs[295]), .I3(
        regs[263]), .S0(n49), .S1(n78), .Z(n580) );
  MUX4V2_8TH40 U616 ( .I0(regs[872]), .I1(regs[840]), .I2(regs[808]), .I3(
        regs[776]), .S0(n50), .S1(n79), .Z(n595) );
  MUX4V2_8TH40 U617 ( .I0(regs[360]), .I1(regs[328]), .I2(regs[296]), .I3(
        regs[264]), .S0(n50), .S1(n78), .Z(n590) );
  MUX4V2_8TH40 U618 ( .I0(regs[873]), .I1(regs[841]), .I2(regs[809]), .I3(
        regs[777]), .S0(n48), .S1(n79), .Z(n605) );
  MUX4V2_8TH40 U619 ( .I0(regs[361]), .I1(regs[329]), .I2(regs[297]), .I3(
        regs[265]), .S0(n50), .S1(n79), .Z(n600) );
  MUX4V2_8TH40 U620 ( .I0(regs[874]), .I1(regs[842]), .I2(regs[810]), .I3(
        regs[778]), .S0(n53), .S1(n80), .Z(n615) );
  MUX4V2_8TH40 U621 ( .I0(regs[362]), .I1(regs[330]), .I2(regs[298]), .I3(
        regs[266]), .S0(n55), .S1(n80), .Z(n610) );
  MUX4V2_8TH40 U622 ( .I0(regs[875]), .I1(regs[843]), .I2(regs[811]), .I3(
        regs[779]), .S0(n56), .S1(n81), .Z(n625) );
  MUX4V2_8TH40 U623 ( .I0(regs[363]), .I1(regs[331]), .I2(regs[299]), .I3(
        regs[267]), .S0(raddr1[0]), .S1(n80), .Z(n620) );
  MUX4V2_8TH40 U624 ( .I0(regs[876]), .I1(regs[844]), .I2(regs[812]), .I3(
        regs[780]), .S0(n56), .S1(n81), .Z(n635) );
  MUX4V2_8TH40 U625 ( .I0(regs[364]), .I1(regs[332]), .I2(regs[300]), .I3(
        regs[268]), .S0(raddr1[0]), .S1(n81), .Z(n630) );
  MUX4V2_8TH40 U626 ( .I0(regs[877]), .I1(regs[845]), .I2(regs[813]), .I3(
        regs[781]), .S0(n51), .S1(n82), .Z(n645) );
  MUX4V2_8TH40 U627 ( .I0(regs[365]), .I1(regs[333]), .I2(regs[301]), .I3(
        regs[269]), .S0(n51), .S1(n81), .Z(n640) );
  MUX4V2_8TH40 U628 ( .I0(regs[878]), .I1(regs[846]), .I2(regs[814]), .I3(
        regs[782]), .S0(n52), .S1(n82), .Z(n655) );
  MUX4V2_8TH40 U629 ( .I0(regs[366]), .I1(regs[334]), .I2(regs[302]), .I3(
        regs[270]), .S0(n51), .S1(n82), .Z(n650) );
  MUX4V2_8TH40 U630 ( .I0(regs[879]), .I1(regs[847]), .I2(regs[815]), .I3(
        regs[783]), .S0(n52), .S1(raddr1[1]), .Z(n665) );
  MUX4V2_8TH40 U631 ( .I0(regs[367]), .I1(regs[335]), .I2(regs[303]), .I3(
        regs[271]), .S0(n52), .S1(raddr1[1]), .Z(n660) );
  MUX4V2_8TH40 U632 ( .I0(regs[368]), .I1(regs[336]), .I2(regs[304]), .I3(
        regs[272]), .S0(n53), .S1(n68), .Z(n670) );
  MUX4V2_8TH40 U633 ( .I0(regs[369]), .I1(regs[337]), .I2(regs[305]), .I3(
        regs[273]), .S0(n53), .S1(n68), .Z(n680) );
  MUX4V2_8TH40 U634 ( .I0(regs[370]), .I1(regs[338]), .I2(regs[306]), .I3(
        regs[274]), .S0(n53), .S1(n69), .Z(n690) );
  MUX4V2_8TH40 U635 ( .I0(regs[371]), .I1(regs[339]), .I2(regs[307]), .I3(
        regs[275]), .S0(raddr1[0]), .S1(n70), .Z(n700) );
  MUX4V2_8TH40 U636 ( .I0(regs[372]), .I1(regs[340]), .I2(regs[308]), .I3(
        regs[276]), .S0(n54), .S1(n70), .Z(n710) );
  MUX4V2_8TH40 U637 ( .I0(regs[373]), .I1(regs[341]), .I2(regs[309]), .I3(
        regs[277]), .S0(n51), .S1(n71), .Z(n720) );
  MUX4V2_8TH40 U638 ( .I0(regs[374]), .I1(regs[342]), .I2(regs[310]), .I3(
        regs[278]), .S0(n52), .S1(n71), .Z(n730) );
  MUX4V2_8TH40 U639 ( .I0(regs[375]), .I1(regs[343]), .I2(regs[311]), .I3(
        regs[279]), .S0(n55), .S1(n76), .Z(n740) );
  MUX4V2_8TH40 U640 ( .I0(regs[376]), .I1(regs[344]), .I2(regs[312]), .I3(
        regs[280]), .S0(n55), .S1(n72), .Z(n750) );
  MUX4V2_8TH40 U641 ( .I0(regs[377]), .I1(regs[345]), .I2(regs[313]), .I3(
        regs[281]), .S0(n56), .S1(n73), .Z(n760) );
  MUX4V2_8TH40 U642 ( .I0(regs[378]), .I1(regs[346]), .I2(regs[314]), .I3(
        regs[282]), .S0(n57), .S1(raddr1[1]), .Z(n770) );
  MUX4V2_8TH40 U643 ( .I0(regs[379]), .I1(regs[347]), .I2(regs[315]), .I3(
        regs[283]), .S0(n57), .S1(n68), .Z(n780) );
  MUX4V2_8TH40 U644 ( .I0(regs[380]), .I1(regs[348]), .I2(regs[316]), .I3(
        regs[284]), .S0(n58), .S1(n74), .Z(n790) );
  MUX4V2_8TH40 U645 ( .I0(regs[381]), .I1(regs[349]), .I2(regs[317]), .I3(
        regs[285]), .S0(n54), .S1(n72), .Z(n800) );
  MUX4V2_8TH40 U646 ( .I0(regs[382]), .I1(regs[350]), .I2(regs[318]), .I3(
        regs[286]), .S0(n53), .S1(n72), .Z(n810) );
  MUX4V2_8TH40 U647 ( .I0(regs[895]), .I1(regs[863]), .I2(regs[831]), .I3(
        regs[799]), .S0(n7), .S1(raddr2[1]), .Z(n1145) );
  MUX4V2_8TH40 U648 ( .I0(regs[383]), .I1(regs[351]), .I2(regs[319]), .I3(
        regs[287]), .S0(n8), .S1(n23), .Z(n1140) );
  MUX4V2_8TH40 U649 ( .I0(regs[383]), .I1(regs[351]), .I2(regs[319]), .I3(
        regs[287]), .S0(raddr1[0]), .S1(n73), .Z(n820) );
  MUX4V2_8TH40 U650 ( .I0(regs[608]), .I1(regs[576]), .I2(regs[544]), .I3(
        regs[512]), .S0(n1), .S1(n27), .Z(n833) );
  MUX4V2_8TH40 U651 ( .I0(regs[609]), .I1(regs[577]), .I2(regs[545]), .I3(
        regs[513]), .S0(n1), .S1(n28), .Z(n843) );
  MUX4V2_8TH40 U652 ( .I0(regs[610]), .I1(regs[578]), .I2(regs[546]), .I3(
        regs[514]), .S0(n2), .S1(n32), .Z(n853) );
  MUX4V2_8TH40 U653 ( .I0(regs[611]), .I1(regs[579]), .I2(regs[547]), .I3(
        regs[515]), .S0(n3), .S1(n25), .Z(n863) );
  MUX4V2_8TH40 U654 ( .I0(regs[612]), .I1(regs[580]), .I2(regs[548]), .I3(
        regs[516]), .S0(n3), .S1(n31), .Z(n873) );
  MUX4V2_8TH40 U655 ( .I0(regs[613]), .I1(regs[581]), .I2(regs[549]), .I3(
        regs[517]), .S0(n4), .S1(n32), .Z(n883) );
  MUX4V2_8TH40 U656 ( .I0(regs[614]), .I1(regs[582]), .I2(regs[550]), .I3(
        regs[518]), .S0(n5), .S1(n32), .Z(n893) );
  MUX4V2_8TH40 U657 ( .I0(regs[615]), .I1(regs[583]), .I2(regs[551]), .I3(
        regs[519]), .S0(n5), .S1(n33), .Z(n903) );
  MUX4V2_8TH40 U658 ( .I0(regs[616]), .I1(regs[584]), .I2(regs[552]), .I3(
        regs[520]), .S0(n6), .S1(n34), .Z(n913) );
  MUX4V2_8TH40 U659 ( .I0(regs[617]), .I1(regs[585]), .I2(regs[553]), .I3(
        regs[521]), .S0(n6), .S1(n34), .Z(n923) );
  MUX4V2_8TH40 U660 ( .I0(regs[618]), .I1(regs[586]), .I2(regs[554]), .I3(
        regs[522]), .S0(n7), .S1(n35), .Z(n933) );
  MUX4V2_8TH40 U661 ( .I0(regs[619]), .I1(regs[587]), .I2(regs[555]), .I3(
        regs[523]), .S0(n8), .S1(n35), .Z(n943) );
  MUX4V2_8TH40 U662 ( .I0(regs[620]), .I1(regs[588]), .I2(regs[556]), .I3(
        regs[524]), .S0(n8), .S1(n36), .Z(n953) );
  MUX4V2_8TH40 U663 ( .I0(regs[621]), .I1(regs[589]), .I2(regs[557]), .I3(
        regs[525]), .S0(n9), .S1(n33), .Z(n963) );
  MUX4V2_8TH40 U664 ( .I0(regs[622]), .I1(regs[590]), .I2(regs[558]), .I3(
        regs[526]), .S0(n9), .S1(n34), .Z(n973) );
  MUX4V2_8TH40 U665 ( .I0(regs[623]), .I1(regs[591]), .I2(regs[559]), .I3(
        regs[527]), .S0(n10), .S1(raddr2[1]), .Z(n983) );
  MUX4V2_8TH40 U666 ( .I0(regs[624]), .I1(regs[592]), .I2(regs[560]), .I3(
        regs[528]), .S0(n11), .S1(n23), .Z(n993) );
  MUX4V2_8TH40 U667 ( .I0(regs[112]), .I1(regs[80]), .I2(regs[48]), .I3(
        regs[16]), .S0(n10), .S1(n27), .Z(n988) );
  MUX4V2_8TH40 U668 ( .I0(regs[625]), .I1(regs[593]), .I2(regs[561]), .I3(
        regs[529]), .S0(n11), .S1(n23), .Z(n1003) );
  MUX4V2_8TH40 U669 ( .I0(regs[113]), .I1(regs[81]), .I2(regs[49]), .I3(
        regs[17]), .S0(n11), .S1(n23), .Z(n998) );
  MUX4V2_8TH40 U670 ( .I0(regs[626]), .I1(regs[594]), .I2(regs[562]), .I3(
        regs[530]), .S0(n12), .S1(n24), .Z(n1013) );
  MUX4V2_8TH40 U671 ( .I0(regs[114]), .I1(regs[82]), .I2(regs[50]), .I3(
        regs[18]), .S0(n12), .S1(n24), .Z(n1008) );
  MUX4V2_8TH40 U672 ( .I0(regs[627]), .I1(regs[595]), .I2(regs[563]), .I3(
        regs[531]), .S0(n3), .S1(n25), .Z(n1023) );
  MUX4V2_8TH40 U673 ( .I0(regs[115]), .I1(regs[83]), .I2(regs[51]), .I3(
        regs[19]), .S0(n12), .S1(n24), .Z(n1018) );
  MUX4V2_8TH40 U674 ( .I0(regs[628]), .I1(regs[596]), .I2(regs[564]), .I3(
        regs[532]), .S0(raddr2[0]), .S1(n25), .Z(n1033) );
  MUX4V2_8TH40 U675 ( .I0(regs[116]), .I1(regs[84]), .I2(regs[52]), .I3(
        regs[20]), .S0(n5), .S1(n25), .Z(n1028) );
  MUX4V2_8TH40 U676 ( .I0(regs[629]), .I1(regs[597]), .I2(regs[565]), .I3(
        regs[533]), .S0(n9), .S1(n26), .Z(n1043) );
  MUX4V2_8TH40 U677 ( .I0(regs[117]), .I1(regs[85]), .I2(regs[53]), .I3(
        regs[21]), .S0(n6), .S1(n26), .Z(n1038) );
  MUX4V2_8TH40 U678 ( .I0(regs[630]), .I1(regs[598]), .I2(regs[566]), .I3(
        regs[534]), .S0(n10), .S1(n27), .Z(n1053) );
  MUX4V2_8TH40 U679 ( .I0(regs[118]), .I1(regs[86]), .I2(regs[54]), .I3(
        regs[22]), .S0(n1), .S1(n26), .Z(n1048) );
  MUX4V2_8TH40 U680 ( .I0(regs[631]), .I1(regs[599]), .I2(regs[567]), .I3(
        regs[535]), .S0(raddr2[0]), .S1(n27), .Z(n1063) );
  MUX4V2_8TH40 U681 ( .I0(regs[119]), .I1(regs[87]), .I2(regs[55]), .I3(
        regs[23]), .S0(n5), .S1(n27), .Z(n1058) );
  MUX4V2_8TH40 U682 ( .I0(regs[632]), .I1(regs[600]), .I2(regs[568]), .I3(
        regs[536]), .S0(n3), .S1(n28), .Z(n1073) );
  MUX4V2_8TH40 U683 ( .I0(regs[120]), .I1(regs[88]), .I2(regs[56]), .I3(
        regs[24]), .S0(n6), .S1(n28), .Z(n1068) );
  MUX4V2_8TH40 U684 ( .I0(regs[633]), .I1(regs[601]), .I2(regs[569]), .I3(
        regs[537]), .S0(raddr2[0]), .S1(n28), .Z(n1083) );
  MUX4V2_8TH40 U685 ( .I0(regs[121]), .I1(regs[89]), .I2(regs[57]), .I3(
        regs[25]), .S0(n5), .S1(n28), .Z(n1078) );
  MUX4V2_8TH40 U686 ( .I0(regs[634]), .I1(regs[602]), .I2(regs[570]), .I3(
        regs[538]), .S0(n13), .S1(n29), .Z(n1093) );
  MUX4V2_8TH40 U687 ( .I0(regs[122]), .I1(regs[90]), .I2(regs[58]), .I3(
        regs[26]), .S0(n13), .S1(n29), .Z(n1088) );
  MUX4V2_8TH40 U688 ( .I0(regs[635]), .I1(regs[603]), .I2(regs[571]), .I3(
        regs[539]), .S0(n13), .S1(n30), .Z(n1103) );
  MUX4V2_8TH40 U689 ( .I0(regs[123]), .I1(regs[91]), .I2(regs[59]), .I3(
        regs[27]), .S0(n13), .S1(n29), .Z(n1098) );
  MUX4V2_8TH40 U690 ( .I0(regs[636]), .I1(regs[604]), .I2(regs[572]), .I3(
        regs[540]), .S0(n14), .S1(n30), .Z(n1113) );
  MUX4V2_8TH40 U691 ( .I0(regs[124]), .I1(regs[92]), .I2(regs[60]), .I3(
        regs[28]), .S0(n14), .S1(n30), .Z(n1108) );
  MUX4V2_8TH40 U692 ( .I0(regs[637]), .I1(regs[605]), .I2(regs[573]), .I3(
        regs[541]), .S0(raddr2[0]), .S1(n23), .Z(n1123) );
  MUX4V2_8TH40 U693 ( .I0(regs[125]), .I1(regs[93]), .I2(regs[61]), .I3(
        regs[29]), .S0(n14), .S1(n24), .Z(n1118) );
  MUX4V2_8TH40 U694 ( .I0(regs[638]), .I1(regs[606]), .I2(regs[574]), .I3(
        regs[542]), .S0(n5), .S1(n27), .Z(n1133) );
  MUX4V2_8TH40 U695 ( .I0(regs[126]), .I1(regs[94]), .I2(regs[62]), .I3(
        regs[30]), .S0(raddr2[0]), .S1(n28), .Z(n1128) );
  MUX4V2_8TH40 U696 ( .I0(regs[608]), .I1(regs[576]), .I2(regs[544]), .I3(
        regs[512]), .S0(n45), .S1(n74), .Z(n97) );
  MUX4V2_8TH40 U697 ( .I0(regs[96]), .I1(regs[64]), .I2(regs[32]), .I3(regs[0]), .S0(n45), .S1(n68), .Z(n92) );
  MUX4V2_8TH40 U698 ( .I0(regs[609]), .I1(regs[577]), .I2(regs[545]), .I3(
        regs[513]), .S0(n45), .S1(n74), .Z(n107) );
  MUX4V2_8TH40 U699 ( .I0(regs[97]), .I1(regs[65]), .I2(regs[33]), .I3(regs[1]), .S0(n45), .S1(n74), .Z(n102) );
  MUX4V2_8TH40 U700 ( .I0(regs[610]), .I1(regs[578]), .I2(regs[546]), .I3(
        regs[514]), .S0(n46), .S1(n75), .Z(n533) );
  MUX4V2_8TH40 U701 ( .I0(regs[98]), .I1(regs[66]), .I2(regs[34]), .I3(regs[2]), .S0(n46), .S1(n75), .Z(n112) );
  MUX4V2_8TH40 U702 ( .I0(regs[611]), .I1(regs[579]), .I2(regs[547]), .I3(
        regs[515]), .S0(n47), .S1(n75), .Z(n543) );
  MUX4V2_8TH40 U703 ( .I0(regs[99]), .I1(regs[67]), .I2(regs[35]), .I3(regs[3]), .S0(n46), .S1(n75), .Z(n538) );
  MUX4V2_8TH40 U704 ( .I0(regs[612]), .I1(regs[580]), .I2(regs[548]), .I3(
        regs[516]), .S0(n47), .S1(n76), .Z(n553) );
  MUX4V2_8TH40 U705 ( .I0(regs[100]), .I1(regs[68]), .I2(regs[36]), .I3(
        regs[4]), .S0(n47), .S1(n76), .Z(n548) );
  MUX4V2_8TH40 U706 ( .I0(regs[613]), .I1(regs[581]), .I2(regs[549]), .I3(
        regs[517]), .S0(n48), .S1(n77), .Z(n563) );
  MUX4V2_8TH40 U707 ( .I0(regs[614]), .I1(regs[582]), .I2(regs[550]), .I3(
        regs[518]), .S0(n49), .S1(n77), .Z(n573) );
  MUX4V2_8TH40 U708 ( .I0(regs[615]), .I1(regs[583]), .I2(regs[551]), .I3(
        regs[519]), .S0(n49), .S1(n78), .Z(n583) );
  MUX4V2_8TH40 U709 ( .I0(regs[616]), .I1(regs[584]), .I2(regs[552]), .I3(
        regs[520]), .S0(n50), .S1(n79), .Z(n593) );
  MUX4V2_8TH40 U710 ( .I0(regs[617]), .I1(regs[585]), .I2(regs[553]), .I3(
        regs[521]), .S0(n50), .S1(n79), .Z(n603) );
  MUX4V2_8TH40 U711 ( .I0(regs[618]), .I1(regs[586]), .I2(regs[554]), .I3(
        regs[522]), .S0(n54), .S1(n80), .Z(n613) );
  MUX4V2_8TH40 U712 ( .I0(regs[619]), .I1(regs[587]), .I2(regs[555]), .I3(
        regs[523]), .S0(n54), .S1(n80), .Z(n623) );
  MUX4V2_8TH40 U713 ( .I0(regs[620]), .I1(regs[588]), .I2(regs[556]), .I3(
        regs[524]), .S0(n55), .S1(n81), .Z(n633) );
  MUX4V2_8TH40 U714 ( .I0(regs[621]), .I1(regs[589]), .I2(regs[557]), .I3(
        regs[525]), .S0(n51), .S1(n82), .Z(n643) );
  MUX4V2_8TH40 U715 ( .I0(regs[622]), .I1(regs[590]), .I2(regs[558]), .I3(
        regs[526]), .S0(n51), .S1(n82), .Z(n653) );
  MUX4V2_8TH40 U716 ( .I0(regs[623]), .I1(regs[591]), .I2(regs[559]), .I3(
        regs[527]), .S0(n52), .S1(raddr1[1]), .Z(n663) );
  MUX4V2_8TH40 U717 ( .I0(regs[112]), .I1(regs[80]), .I2(regs[48]), .I3(
        regs[16]), .S0(n52), .S1(n77), .Z(n668) );
  MUX4V2_8TH40 U718 ( .I0(regs[113]), .I1(regs[81]), .I2(regs[49]), .I3(
        regs[17]), .S0(n53), .S1(n68), .Z(n678) );
  MUX4V2_8TH40 U719 ( .I0(regs[114]), .I1(regs[82]), .I2(regs[50]), .I3(
        regs[18]), .S0(n54), .S1(n69), .Z(n688) );
  MUX4V2_8TH40 U720 ( .I0(regs[115]), .I1(regs[83]), .I2(regs[51]), .I3(
        regs[19]), .S0(n55), .S1(n69), .Z(n698) );
  MUX4V2_8TH40 U721 ( .I0(regs[116]), .I1(regs[84]), .I2(regs[52]), .I3(
        regs[20]), .S0(n54), .S1(n70), .Z(n708) );
  MUX4V2_8TH40 U722 ( .I0(regs[117]), .I1(regs[85]), .I2(regs[53]), .I3(
        regs[21]), .S0(n54), .S1(n71), .Z(n718) );
  MUX4V2_8TH40 U723 ( .I0(regs[118]), .I1(regs[86]), .I2(regs[54]), .I3(
        regs[22]), .S0(n45), .S1(n71), .Z(n728) );
  MUX4V2_8TH40 U724 ( .I0(regs[119]), .I1(regs[87]), .I2(regs[55]), .I3(
        regs[23]), .S0(n55), .S1(n70), .Z(n738) );
  MUX4V2_8TH40 U725 ( .I0(regs[120]), .I1(regs[88]), .I2(regs[56]), .I3(
        regs[24]), .S0(n55), .S1(n78), .Z(n748) );
  MUX4V2_8TH40 U726 ( .I0(regs[121]), .I1(regs[89]), .I2(regs[57]), .I3(
        regs[25]), .S0(n56), .S1(n79), .Z(n758) );
  MUX4V2_8TH40 U727 ( .I0(regs[122]), .I1(regs[90]), .I2(regs[58]), .I3(
        regs[26]), .S0(n57), .S1(n69), .Z(n768) );
  MUX4V2_8TH40 U728 ( .I0(regs[123]), .I1(regs[91]), .I2(regs[59]), .I3(
        regs[27]), .S0(n57), .S1(n74), .Z(n778) );
  MUX4V2_8TH40 U729 ( .I0(regs[124]), .I1(regs[92]), .I2(regs[60]), .I3(
        regs[28]), .S0(n58), .S1(n75), .Z(n788) );
  MUX4V2_8TH40 U730 ( .I0(regs[125]), .I1(regs[93]), .I2(regs[61]), .I3(
        regs[29]), .S0(n58), .S1(n72), .Z(n798) );
  MUX4V2_8TH40 U731 ( .I0(regs[126]), .I1(regs[94]), .I2(regs[62]), .I3(
        regs[30]), .S0(n57), .S1(n72), .Z(n808) );
  MUX4V2_8TH40 U732 ( .I0(regs[639]), .I1(regs[607]), .I2(regs[575]), .I3(
        regs[543]), .S0(n11), .S1(n24), .Z(n1143) );
  MUX4V2_8TH40 U733 ( .I0(regs[127]), .I1(regs[95]), .I2(regs[63]), .I3(
        regs[31]), .S0(n12), .S1(n27), .Z(n1138) );
  MUX4V2_8TH40 U734 ( .I0(regs[127]), .I1(regs[95]), .I2(regs[63]), .I3(
        regs[31]), .S0(raddr1[0]), .S1(n73), .Z(n818) );
  MUX4V4_8TH40 U735 ( .I0(n95), .I1(n93), .I2(n94), .I3(n92), .S0(raddr1[3]), 
        .S1(raddr1[2]), .Z(n96) );
  MUX4V4_8TH40 U736 ( .I0(n100), .I1(n98), .I2(n99), .I3(n97), .S0(raddr1[3]), 
        .S1(raddr1[2]), .Z(n101) );
  MUX4V4_8TH40 U737 ( .I0(n105), .I1(n103), .I2(n104), .I3(n102), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n106) );
  MUX4V4_8TH40 U738 ( .I0(n110), .I1(n108), .I2(n109), .I3(n107), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n111) );
  MUX4V4_8TH40 U739 ( .I0(n531), .I1(n529), .I2(n530), .I3(n112), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n532) );
  MUX4V4_8TH40 U740 ( .I0(n536), .I1(n534), .I2(n535), .I3(n533), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n537) );
  MUX4V4_8TH40 U741 ( .I0(n541), .I1(n539), .I2(n540), .I3(n538), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n542) );
  MUX4V4_8TH40 U742 ( .I0(n546), .I1(n544), .I2(n545), .I3(n543), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n547) );
  MUX4V4_8TH40 U743 ( .I0(n551), .I1(n549), .I2(n550), .I3(n548), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n552) );
  MUX4V4_8TH40 U744 ( .I0(n556), .I1(n554), .I2(n555), .I3(n553), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n557) );
  MUX4V4_8TH40 U745 ( .I0(n561), .I1(n559), .I2(n560), .I3(n558), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n562) );
  MUX4V4_8TH40 U746 ( .I0(n566), .I1(n564), .I2(n565), .I3(n563), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n567) );
  MUX4V4_8TH40 U747 ( .I0(n571), .I1(n569), .I2(n570), .I3(n568), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n572) );
  MUX4V4_8TH40 U748 ( .I0(n576), .I1(n574), .I2(n575), .I3(n573), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n577) );
  MUX4V4_8TH40 U749 ( .I0(n581), .I1(n579), .I2(n580), .I3(n578), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n582) );
  MUX4V4_8TH40 U750 ( .I0(n586), .I1(n584), .I2(n585), .I3(n583), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n587) );
  MUX4V4_8TH40 U751 ( .I0(n591), .I1(n589), .I2(n590), .I3(n588), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n592) );
  MUX4V4_8TH40 U752 ( .I0(n596), .I1(n594), .I2(n595), .I3(n593), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n597) );
  MUX4V4_8TH40 U753 ( .I0(n601), .I1(n599), .I2(n600), .I3(n598), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n602) );
  MUX4V4_8TH40 U754 ( .I0(n606), .I1(n604), .I2(n605), .I3(n603), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n607) );
  MUX4V4_8TH40 U755 ( .I0(n611), .I1(n609), .I2(n610), .I3(n608), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n612) );
  MUX4V4_8TH40 U756 ( .I0(n616), .I1(n614), .I2(n615), .I3(n613), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n617) );
  MUX4V4_8TH40 U757 ( .I0(n621), .I1(n619), .I2(n620), .I3(n618), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n622) );
  MUX4V4_8TH40 U758 ( .I0(n626), .I1(n624), .I2(n625), .I3(n623), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n627) );
  MUX4V4_8TH40 U759 ( .I0(n631), .I1(n629), .I2(n630), .I3(n628), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n632) );
  MUX4V4_8TH40 U760 ( .I0(n636), .I1(n634), .I2(n635), .I3(n633), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n637) );
  MUX4V4_8TH40 U761 ( .I0(n641), .I1(n639), .I2(n640), .I3(n638), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n642) );
  MUX4V4_8TH40 U762 ( .I0(n646), .I1(n644), .I2(n645), .I3(n643), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n647) );
  MUX4V4_8TH40 U763 ( .I0(n651), .I1(n649), .I2(n650), .I3(n648), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n652) );
  MUX4V4_8TH40 U764 ( .I0(n656), .I1(n654), .I2(n655), .I3(n653), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n657) );
  MUX4V4_8TH40 U765 ( .I0(n661), .I1(n659), .I2(n660), .I3(n658), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n662) );
  MUX4V4_8TH40 U766 ( .I0(n666), .I1(n664), .I2(n665), .I3(n663), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n667) );
  MUX4V4_8TH40 U767 ( .I0(n671), .I1(n669), .I2(n670), .I3(n668), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n672) );
  MUX4V4_8TH40 U768 ( .I0(n676), .I1(n674), .I2(n675), .I3(n673), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n677) );
  CKMUX2V4_8TH40 U769 ( .I0(n677), .I1(n672), .S(raddr1[4]), .Z(N110) );
  MUX4V4_8TH40 U770 ( .I0(n681), .I1(n679), .I2(n680), .I3(n678), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n682) );
  MUX4V4_8TH40 U771 ( .I0(n686), .I1(n684), .I2(n685), .I3(n683), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n687) );
  CKMUX2V4_8TH40 U772 ( .I0(n687), .I1(n682), .S(raddr1[4]), .Z(N109) );
  MUX4V4_8TH40 U773 ( .I0(n691), .I1(n689), .I2(n690), .I3(n688), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n692) );
  MUX4V4_8TH40 U774 ( .I0(n696), .I1(n694), .I2(n695), .I3(n693), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n697) );
  CKMUX2V4_8TH40 U775 ( .I0(n697), .I1(n692), .S(raddr1[4]), .Z(N108) );
  MUX4V4_8TH40 U776 ( .I0(n701), .I1(n699), .I2(n700), .I3(n698), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n702) );
  MUX4V4_8TH40 U777 ( .I0(n706), .I1(n704), .I2(n705), .I3(n703), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n707) );
  CKMUX2V4_8TH40 U778 ( .I0(n707), .I1(n702), .S(raddr1[4]), .Z(N107) );
  MUX4V4_8TH40 U779 ( .I0(n711), .I1(n709), .I2(n710), .I3(n708), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n712) );
  MUX4V4_8TH40 U780 ( .I0(n716), .I1(n714), .I2(n715), .I3(n713), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n717) );
  CKMUX2V4_8TH40 U781 ( .I0(n717), .I1(n712), .S(raddr1[4]), .Z(N106) );
  MUX4V4_8TH40 U782 ( .I0(n721), .I1(n719), .I2(n720), .I3(n718), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n722) );
  MUX4V4_8TH40 U783 ( .I0(n726), .I1(n724), .I2(n725), .I3(n723), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n727) );
  CKMUX2V4_8TH40 U784 ( .I0(n727), .I1(n722), .S(raddr1[4]), .Z(N105) );
  MUX4V4_8TH40 U785 ( .I0(n731), .I1(n729), .I2(n730), .I3(n728), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n732) );
  MUX4V4_8TH40 U786 ( .I0(n736), .I1(n734), .I2(n735), .I3(n733), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n737) );
  CKMUX2V4_8TH40 U787 ( .I0(n737), .I1(n732), .S(raddr1[4]), .Z(N104) );
  MUX4V4_8TH40 U788 ( .I0(n741), .I1(n739), .I2(n740), .I3(n738), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n742) );
  MUX4V4_8TH40 U789 ( .I0(n746), .I1(n744), .I2(n745), .I3(n743), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n747) );
  CKMUX2V4_8TH40 U790 ( .I0(n747), .I1(n742), .S(raddr1[4]), .Z(N103) );
  MUX4V4_8TH40 U791 ( .I0(n751), .I1(n749), .I2(n750), .I3(n748), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n752) );
  MUX4V4_8TH40 U792 ( .I0(n756), .I1(n754), .I2(n755), .I3(n753), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n757) );
  CKMUX2V4_8TH40 U793 ( .I0(n757), .I1(n752), .S(raddr1[4]), .Z(N102) );
  MUX4V4_8TH40 U794 ( .I0(n761), .I1(n759), .I2(n760), .I3(n758), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n762) );
  MUX4V4_8TH40 U795 ( .I0(n766), .I1(n764), .I2(n765), .I3(n763), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n767) );
  CKMUX2V4_8TH40 U796 ( .I0(n767), .I1(n762), .S(raddr1[4]), .Z(N101) );
  MUX4V4_8TH40 U797 ( .I0(n771), .I1(n769), .I2(n770), .I3(n768), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n772) );
  MUX4V4_8TH40 U798 ( .I0(n776), .I1(n774), .I2(n775), .I3(n773), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n777) );
  CKMUX2V4_8TH40 U799 ( .I0(n777), .I1(n772), .S(raddr1[4]), .Z(N100) );
  MUX4V4_8TH40 U800 ( .I0(n781), .I1(n779), .I2(n780), .I3(n778), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n782) );
  MUX4V4_8TH40 U801 ( .I0(n786), .I1(n784), .I2(n785), .I3(n783), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n787) );
  CKMUX2V4_8TH40 U802 ( .I0(n787), .I1(n782), .S(raddr1[4]), .Z(N99) );
  MUX4V4_8TH40 U803 ( .I0(n791), .I1(n789), .I2(n790), .I3(n788), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n792) );
  MUX4V4_8TH40 U804 ( .I0(n796), .I1(n794), .I2(n795), .I3(n793), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n797) );
  CKMUX2V4_8TH40 U805 ( .I0(n797), .I1(n792), .S(raddr1[4]), .Z(N98) );
  MUX4V4_8TH40 U806 ( .I0(n801), .I1(n799), .I2(n800), .I3(n798), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n802) );
  MUX4V4_8TH40 U807 ( .I0(n806), .I1(n804), .I2(n805), .I3(n803), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n807) );
  CKMUX2V4_8TH40 U808 ( .I0(n807), .I1(n802), .S(raddr1[4]), .Z(N97) );
  MUX4V4_8TH40 U809 ( .I0(n811), .I1(n809), .I2(n810), .I3(n808), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n812) );
  MUX4V4_8TH40 U810 ( .I0(n816), .I1(n814), .I2(n815), .I3(n813), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n817) );
  CKMUX2V4_8TH40 U811 ( .I0(n817), .I1(n812), .S(raddr1[4]), .Z(N96) );
  MUX4V4_8TH40 U812 ( .I0(n821), .I1(n819), .I2(n820), .I3(n818), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n822) );
  MUX4V4_8TH40 U813 ( .I0(n826), .I1(n824), .I2(n825), .I3(n823), .S0(
        raddr1[3]), .S1(raddr1[2]), .Z(n827) );
  CKMUX2V4_8TH40 U814 ( .I0(n827), .I1(n822), .S(raddr1[4]), .Z(N95) );
  MUX4V4_8TH40 U815 ( .I0(n831), .I1(n829), .I2(n830), .I3(n828), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n832) );
  MUX4V4_8TH40 U816 ( .I0(n836), .I1(n834), .I2(n835), .I3(n833), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n837) );
  MUX4V4_8TH40 U817 ( .I0(n841), .I1(n839), .I2(n840), .I3(n838), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n842) );
  MUX4V4_8TH40 U818 ( .I0(n846), .I1(n844), .I2(n845), .I3(n843), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n847) );
  MUX4V4_8TH40 U819 ( .I0(n851), .I1(n849), .I2(n850), .I3(n848), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n852) );
  MUX4V4_8TH40 U820 ( .I0(n856), .I1(n854), .I2(n855), .I3(n853), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n857) );
  MUX4V4_8TH40 U821 ( .I0(n861), .I1(n859), .I2(n860), .I3(n858), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n862) );
  MUX4V4_8TH40 U822 ( .I0(n866), .I1(n864), .I2(n865), .I3(n863), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n867) );
  MUX4V4_8TH40 U823 ( .I0(n871), .I1(n869), .I2(n870), .I3(n868), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n872) );
  MUX4V4_8TH40 U824 ( .I0(n876), .I1(n874), .I2(n875), .I3(n873), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n877) );
  MUX4V4_8TH40 U825 ( .I0(n881), .I1(n879), .I2(n880), .I3(n878), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n882) );
  MUX4V4_8TH40 U826 ( .I0(n886), .I1(n884), .I2(n885), .I3(n883), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n887) );
  MUX4V4_8TH40 U827 ( .I0(n891), .I1(n889), .I2(n890), .I3(n888), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n892) );
  MUX4V4_8TH40 U828 ( .I0(n896), .I1(n894), .I2(n895), .I3(n893), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n897) );
  MUX4V4_8TH40 U829 ( .I0(n901), .I1(n899), .I2(n900), .I3(n898), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n902) );
  MUX4V4_8TH40 U830 ( .I0(n906), .I1(n904), .I2(n905), .I3(n903), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n907) );
  MUX4V4_8TH40 U831 ( .I0(n911), .I1(n909), .I2(n910), .I3(n908), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n912) );
  MUX4V4_8TH40 U832 ( .I0(n916), .I1(n914), .I2(n915), .I3(n913), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n917) );
  MUX4V4_8TH40 U833 ( .I0(n921), .I1(n919), .I2(n920), .I3(n918), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n922) );
  MUX4V4_8TH40 U834 ( .I0(n926), .I1(n924), .I2(n925), .I3(n923), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n927) );
  MUX4V4_8TH40 U835 ( .I0(n931), .I1(n929), .I2(n930), .I3(n928), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n932) );
  MUX4V4_8TH40 U836 ( .I0(n936), .I1(n934), .I2(n935), .I3(n933), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n937) );
  MUX4V4_8TH40 U837 ( .I0(n941), .I1(n939), .I2(n940), .I3(n938), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n942) );
  MUX4V4_8TH40 U838 ( .I0(n946), .I1(n944), .I2(n945), .I3(n943), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n947) );
  MUX4V4_8TH40 U839 ( .I0(n951), .I1(n949), .I2(n950), .I3(n948), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n952) );
  MUX4V4_8TH40 U840 ( .I0(n956), .I1(n954), .I2(n955), .I3(n953), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n957) );
  MUX4V4_8TH40 U841 ( .I0(n961), .I1(n959), .I2(n960), .I3(n958), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n962) );
  MUX4V4_8TH40 U842 ( .I0(n966), .I1(n964), .I2(n965), .I3(n963), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n967) );
  MUX4V4_8TH40 U843 ( .I0(n971), .I1(n969), .I2(n970), .I3(n968), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n972) );
  MUX4V4_8TH40 U844 ( .I0(n976), .I1(n974), .I2(n975), .I3(n973), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n977) );
  MUX4V4_8TH40 U845 ( .I0(n981), .I1(n979), .I2(n980), .I3(n978), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n982) );
  MUX4V4_8TH40 U846 ( .I0(n986), .I1(n984), .I2(n985), .I3(n983), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n987) );
  MUX4V4_8TH40 U847 ( .I0(n991), .I1(n989), .I2(n990), .I3(n988), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n992) );
  MUX4V4_8TH40 U848 ( .I0(n996), .I1(n994), .I2(n995), .I3(n993), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n997) );
  MUX4V4_8TH40 U849 ( .I0(n1001), .I1(n999), .I2(n1000), .I3(n998), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1002) );
  MUX4V4_8TH40 U850 ( .I0(n1006), .I1(n1004), .I2(n1005), .I3(n1003), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1007) );
  MUX4V4_8TH40 U851 ( .I0(n1011), .I1(n1009), .I2(n1010), .I3(n1008), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1012) );
  MUX4V4_8TH40 U852 ( .I0(n1016), .I1(n1014), .I2(n1015), .I3(n1013), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1017) );
  MUX4V4_8TH40 U853 ( .I0(n1021), .I1(n1019), .I2(n1020), .I3(n1018), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1022) );
  MUX4V4_8TH40 U854 ( .I0(n1026), .I1(n1024), .I2(n1025), .I3(n1023), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1027) );
  MUX4V4_8TH40 U855 ( .I0(n1031), .I1(n1029), .I2(n1030), .I3(n1028), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1032) );
  MUX4V4_8TH40 U856 ( .I0(n1036), .I1(n1034), .I2(n1035), .I3(n1033), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1037) );
  MUX4V4_8TH40 U857 ( .I0(n1041), .I1(n1039), .I2(n1040), .I3(n1038), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1042) );
  MUX4V4_8TH40 U858 ( .I0(n1046), .I1(n1044), .I2(n1045), .I3(n1043), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1047) );
  MUX4V4_8TH40 U859 ( .I0(n1051), .I1(n1049), .I2(n1050), .I3(n1048), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1052) );
  MUX4V4_8TH40 U860 ( .I0(n1056), .I1(n1054), .I2(n1055), .I3(n1053), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1057) );
  MUX4V4_8TH40 U861 ( .I0(n1061), .I1(n1059), .I2(n1060), .I3(n1058), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1062) );
  MUX4V4_8TH40 U862 ( .I0(n1066), .I1(n1064), .I2(n1065), .I3(n1063), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1067) );
  MUX4V4_8TH40 U863 ( .I0(n1071), .I1(n1069), .I2(n1070), .I3(n1068), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1072) );
  MUX4V4_8TH40 U864 ( .I0(n1076), .I1(n1074), .I2(n1075), .I3(n1073), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1077) );
  MUX4V4_8TH40 U865 ( .I0(n1081), .I1(n1079), .I2(n1080), .I3(n1078), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1082) );
  MUX4V4_8TH40 U866 ( .I0(n1086), .I1(n1084), .I2(n1085), .I3(n1083), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1087) );
  MUX4V4_8TH40 U867 ( .I0(n1091), .I1(n1089), .I2(n1090), .I3(n1088), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1092) );
  MUX4V4_8TH40 U868 ( .I0(n1096), .I1(n1094), .I2(n1095), .I3(n1093), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1097) );
  MUX4V4_8TH40 U869 ( .I0(n1101), .I1(n1099), .I2(n1100), .I3(n1098), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1102) );
  MUX4V4_8TH40 U870 ( .I0(n1106), .I1(n1104), .I2(n1105), .I3(n1103), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1107) );
  MUX4V4_8TH40 U871 ( .I0(n1111), .I1(n1109), .I2(n1110), .I3(n1108), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1112) );
  MUX4V4_8TH40 U872 ( .I0(n1116), .I1(n1114), .I2(n1115), .I3(n1113), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1117) );
  MUX4V4_8TH40 U873 ( .I0(n1121), .I1(n1119), .I2(n1120), .I3(n1118), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1122) );
  MUX4V4_8TH40 U874 ( .I0(n1126), .I1(n1124), .I2(n1125), .I3(n1123), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1127) );
  MUX4V4_8TH40 U875 ( .I0(n1131), .I1(n1129), .I2(n1130), .I3(n1128), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1132) );
  MUX4V4_8TH40 U876 ( .I0(n1136), .I1(n1134), .I2(n1135), .I3(n1133), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1137) );
  MUX4V4_8TH40 U877 ( .I0(n1141), .I1(n1139), .I2(n1140), .I3(n1138), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1142) );
  MUX4V4_8TH40 U878 ( .I0(n1146), .I1(n1144), .I2(n1145), .I3(n1143), .S0(
        raddr2[3]), .S1(raddr2[2]), .Z(n1147) );
  IOA22V0_8TH40 U879 ( .B1(n1148), .B2(n1157), .A1(N140), .A2(n1150), .ZN(
        rdata2[31]) );
  IOA22V0_8TH40 U880 ( .B1(n1148), .B2(n1158), .A1(N141), .A2(n1150), .ZN(
        rdata2[30]) );
  IOA22V0_8TH40 U881 ( .B1(n1148), .B2(n1160), .A1(N142), .A2(n1150), .ZN(
        rdata2[29]) );
  IOA22V0_8TH40 U882 ( .B1(n1148), .B2(n1161), .A1(N143), .A2(n1150), .ZN(
        rdata2[28]) );
  IOA22V0_8TH40 U883 ( .B1(n1148), .B2(n1162), .A1(N144), .A2(n1150), .ZN(
        rdata2[27]) );
  IOA22V0_8TH40 U884 ( .B1(n1148), .B2(n1163), .A1(N145), .A2(n1150), .ZN(
        rdata2[26]) );
  IOA22V0_8TH40 U885 ( .B1(n1148), .B2(n1164), .A1(N146), .A2(n1150), .ZN(
        rdata2[25]) );
  IOA22V0_8TH40 U886 ( .B1(n1148), .B2(n1165), .A1(N147), .A2(n1150), .ZN(
        rdata2[24]) );
  IOA22V0_8TH40 U887 ( .B1(n1148), .B2(n1166), .A1(N148), .A2(n1150), .ZN(
        rdata2[23]) );
  IOA22V0_8TH40 U888 ( .B1(n1148), .B2(n1167), .A1(N149), .A2(n1150), .ZN(
        rdata2[22]) );
  IOA22V0_8TH40 U889 ( .B1(n1148), .B2(n1168), .A1(N150), .A2(n1150), .ZN(
        rdata2[21]) );
  IOA22V0_8TH40 U890 ( .B1(n1148), .B2(n1169), .A1(N151), .A2(n1150), .ZN(
        rdata2[20]) );
  IOA22V0_8TH40 U891 ( .B1(n1148), .B2(n1171), .A1(N152), .A2(n1150), .ZN(
        rdata2[19]) );
  IOA22V0_8TH40 U892 ( .B1(n1148), .B2(n1172), .A1(N153), .A2(n1150), .ZN(
        rdata2[18]) );
  IOA22V0_8TH40 U893 ( .B1(n1148), .B2(n1173), .A1(N154), .A2(n1150), .ZN(
        rdata2[17]) );
  IOA22V0_8TH40 U894 ( .B1(n1148), .B2(n1174), .A1(N155), .A2(n1150), .ZN(
        rdata2[16]) );
  I2NOR4V0_8TH40 U895 ( .A1(re2), .A2(n1182), .B1(n1183), .B2(rst), .ZN(n1150)
         );
  OR3V0_8TH40 U896 ( .A1(n1182), .A2(n1183), .A3(rst), .Z(n1148) );
  XNOR2V0_8TH40 U897 ( .A1(n1191), .A2(raddr2[1]), .ZN(n1190) );
  XNOR2V0_8TH40 U898 ( .A1(n1192), .A2(n4), .ZN(n1189) );
  XNOR2V0_8TH40 U899 ( .A1(raddr2[3]), .A2(waddr[3]), .ZN(n1187) );
  XNOR2V0_8TH40 U900 ( .A1(raddr2[4]), .A2(waddr[4]), .ZN(n1186) );
  XNOR2V0_8TH40 U901 ( .A1(raddr2[2]), .A2(waddr[2]), .ZN(n1185) );
  CLKNV1_8TH40 U902 ( .I(wdata[9]), .ZN(n1149) );
  CLKNV1_8TH40 U903 ( .I(wdata[8]), .ZN(n1151) );
  CLKNV1_8TH40 U904 ( .I(wdata[7]), .ZN(n1152) );
  CLKNV1_8TH40 U905 ( .I(wdata[6]), .ZN(n1153) );
  CLKNV1_8TH40 U906 ( .I(wdata[5]), .ZN(n1154) );
  IOA22V0_8TH40 U907 ( .B1(n1155), .B2(n1193), .A1(N122), .A2(n1194), .ZN(
        rdata1[4]) );
  CLKNV1_8TH40 U908 ( .I(wdata[4]), .ZN(n1155) );
  IOA22V0_8TH40 U909 ( .B1(n1156), .B2(n1193), .A1(N123), .A2(n1194), .ZN(
        rdata1[3]) );
  CLKNV1_8TH40 U910 ( .I(wdata[3]), .ZN(n1156) );
  CLKNV1_8TH40 U911 ( .I(wdata[31]), .ZN(n1157) );
  CLKNV1_8TH40 U912 ( .I(wdata[30]), .ZN(n1158) );
  IOA22V0_8TH40 U913 ( .B1(n1159), .B2(n1193), .A1(N124), .A2(n1194), .ZN(
        rdata1[2]) );
  CLKNV1_8TH40 U914 ( .I(wdata[2]), .ZN(n1159) );
  CLKNV1_8TH40 U915 ( .I(wdata[29]), .ZN(n1160) );
  CLKNV1_8TH40 U916 ( .I(wdata[28]), .ZN(n1161) );
  CLKNV1_8TH40 U917 ( .I(wdata[27]), .ZN(n1162) );
  CLKNV1_8TH40 U918 ( .I(wdata[26]), .ZN(n1163) );
  CLKNV1_8TH40 U919 ( .I(wdata[25]), .ZN(n1164) );
  CLKNV1_8TH40 U920 ( .I(wdata[24]), .ZN(n1165) );
  CLKNV1_8TH40 U921 ( .I(wdata[23]), .ZN(n1166) );
  CLKNV1_8TH40 U922 ( .I(wdata[22]), .ZN(n1167) );
  CLKNV1_8TH40 U923 ( .I(wdata[21]), .ZN(n1168) );
  CLKNV1_8TH40 U924 ( .I(wdata[20]), .ZN(n1169) );
  IOA22V0_8TH40 U925 ( .B1(n1170), .B2(n1193), .A1(N125), .A2(n1194), .ZN(
        rdata1[1]) );
  CLKNV1_8TH40 U926 ( .I(wdata[1]), .ZN(n1170) );
  CLKNV1_8TH40 U927 ( .I(wdata[19]), .ZN(n1171) );
  CLKNV1_8TH40 U928 ( .I(wdata[18]), .ZN(n1172) );
  CLKNV1_8TH40 U929 ( .I(wdata[17]), .ZN(n1173) );
  CLKNV1_8TH40 U930 ( .I(wdata[16]), .ZN(n1174) );
  CLKNV1_8TH40 U931 ( .I(wdata[15]), .ZN(n1175) );
  CLKNV1_8TH40 U932 ( .I(wdata[14]), .ZN(n1176) );
  CLKNV1_8TH40 U933 ( .I(wdata[13]), .ZN(n1177) );
  CLKNV1_8TH40 U934 ( .I(wdata[12]), .ZN(n1178) );
  CLKNV1_8TH40 U935 ( .I(wdata[11]), .ZN(n1179) );
  CLKNV1_8TH40 U936 ( .I(wdata[10]), .ZN(n1180) );
  IOA22V0_8TH40 U937 ( .B1(n1181), .B2(n1193), .A1(N126), .A2(n1194), .ZN(
        rdata1[0]) );
  OR3V0_8TH40 U938 ( .A1(n1195), .A2(n1196), .A3(rst), .Z(n1193) );
  INOR4V0_8TH40 U939 ( .A1(n1197), .B1(raddr1[0]), .B2(raddr1[1]), .B3(
        raddr1[2]), .ZN(n1196) );
  XNOR2V0_8TH40 U940 ( .A1(n1191), .A2(raddr1[1]), .ZN(n1203) );
  XNOR2V0_8TH40 U941 ( .A1(n1192), .A2(raddr1[0]), .ZN(n1202) );
  XNOR2V0_8TH40 U942 ( .A1(raddr1[3]), .A2(waddr[3]), .ZN(n1200) );
  XNOR2V0_8TH40 U943 ( .A1(raddr1[4]), .A2(waddr[4]), .ZN(n1199) );
  XNOR2V0_8TH40 U944 ( .A1(raddr1[2]), .A2(waddr[2]), .ZN(n1198) );
  CLKNV1_8TH40 U945 ( .I(wdata[0]), .ZN(n1181) );
  NAND3V0P5_8TH40 U946 ( .A1(n1191), .A2(n1215), .A3(n1192), .ZN(n1209) );
  NAND3V0P5_8TH40 U947 ( .A1(n1191), .A2(n1215), .A3(waddr[0]), .ZN(n1204) );
  NAND3V0P5_8TH40 U948 ( .A1(n1192), .A2(n1215), .A3(waddr[1]), .ZN(n1206) );
  NAND3V0P5_8TH40 U949 ( .A1(n1192), .A2(n1191), .A3(waddr[2]), .ZN(n1207) );
  CKMUX2V2_8TH40 U950 ( .I0(regs[927]), .I1(wdata[31]), .S(n1216), .Z(n528) );
  CKMUX2V2_8TH40 U951 ( .I0(regs[926]), .I1(wdata[30]), .S(n1216), .Z(n527) );
  CKMUX2V2_8TH40 U952 ( .I0(regs[925]), .I1(wdata[29]), .S(n1216), .Z(n526) );
  CKMUX2V2_8TH40 U953 ( .I0(regs[924]), .I1(wdata[28]), .S(n1216), .Z(n525) );
  CKMUX2V2_8TH40 U954 ( .I0(regs[923]), .I1(wdata[27]), .S(n1216), .Z(n524) );
  CKMUX2V2_8TH40 U955 ( .I0(regs[922]), .I1(wdata[26]), .S(n1216), .Z(n523) );
  CKMUX2V2_8TH40 U956 ( .I0(regs[921]), .I1(wdata[25]), .S(n1216), .Z(n522) );
  CKMUX2V2_8TH40 U957 ( .I0(regs[920]), .I1(wdata[24]), .S(n1216), .Z(n521) );
  CKMUX2V2_8TH40 U958 ( .I0(regs[919]), .I1(wdata[23]), .S(n1216), .Z(n520) );
  CKMUX2V2_8TH40 U959 ( .I0(regs[918]), .I1(wdata[22]), .S(n1216), .Z(n519) );
  CKMUX2V2_8TH40 U960 ( .I0(regs[917]), .I1(wdata[21]), .S(n1216), .Z(n518) );
  CKMUX2V2_8TH40 U961 ( .I0(regs[916]), .I1(wdata[20]), .S(n1216), .Z(n517) );
  CKMUX2V2_8TH40 U962 ( .I0(regs[915]), .I1(wdata[19]), .S(n1216), .Z(n516) );
  CKMUX2V2_8TH40 U963 ( .I0(regs[914]), .I1(wdata[18]), .S(n1216), .Z(n515) );
  CKMUX2V2_8TH40 U964 ( .I0(regs[913]), .I1(wdata[17]), .S(n1216), .Z(n514) );
  CKMUX2V2_8TH40 U965 ( .I0(regs[912]), .I1(wdata[16]), .S(n1216), .Z(n513) );
  CKMUX2V2_8TH40 U966 ( .I0(regs[911]), .I1(wdata[15]), .S(n1216), .Z(n512) );
  CKMUX2V2_8TH40 U967 ( .I0(regs[910]), .I1(wdata[14]), .S(n1216), .Z(n511) );
  CKMUX2V2_8TH40 U968 ( .I0(regs[909]), .I1(wdata[13]), .S(n1216), .Z(n510) );
  CKMUX2V2_8TH40 U969 ( .I0(regs[908]), .I1(wdata[12]), .S(n1216), .Z(n509) );
  CKMUX2V2_8TH40 U970 ( .I0(regs[907]), .I1(wdata[11]), .S(n1216), .Z(n508) );
  CKMUX2V2_8TH40 U971 ( .I0(regs[906]), .I1(wdata[10]), .S(n1216), .Z(n507) );
  CKMUX2V2_8TH40 U972 ( .I0(regs[905]), .I1(wdata[9]), .S(n1216), .Z(n506) );
  CKMUX2V2_8TH40 U973 ( .I0(regs[904]), .I1(wdata[8]), .S(n1216), .Z(n505) );
  CKMUX2V2_8TH40 U974 ( .I0(regs[903]), .I1(wdata[7]), .S(n1216), .Z(n504) );
  CKMUX2V2_8TH40 U975 ( .I0(regs[902]), .I1(wdata[6]), .S(n1216), .Z(n503) );
  CKMUX2V2_8TH40 U976 ( .I0(regs[901]), .I1(wdata[5]), .S(n1216), .Z(n502) );
  CKMUX2V2_8TH40 U977 ( .I0(regs[900]), .I1(wdata[4]), .S(n1216), .Z(n501) );
  CKMUX2V2_8TH40 U978 ( .I0(regs[899]), .I1(wdata[3]), .S(n1216), .Z(n500) );
  CKMUX2V2_8TH40 U979 ( .I0(regs[898]), .I1(wdata[2]), .S(n1216), .Z(n499) );
  CKMUX2V2_8TH40 U980 ( .I0(regs[897]), .I1(wdata[1]), .S(n1216), .Z(n498) );
  CKMUX2V2_8TH40 U981 ( .I0(regs[896]), .I1(wdata[0]), .S(n1216), .Z(n497) );
  CKMUX2V2_8TH40 U982 ( .I0(regs[863]), .I1(wdata[31]), .S(n1217), .Z(n496) );
  CKMUX2V2_8TH40 U983 ( .I0(regs[862]), .I1(wdata[30]), .S(n1217), .Z(n495) );
  CKMUX2V2_8TH40 U984 ( .I0(regs[861]), .I1(wdata[29]), .S(n1217), .Z(n494) );
  CKMUX2V2_8TH40 U985 ( .I0(regs[860]), .I1(wdata[28]), .S(n1217), .Z(n493) );
  CKMUX2V2_8TH40 U986 ( .I0(regs[859]), .I1(wdata[27]), .S(n1217), .Z(n492) );
  CKMUX2V2_8TH40 U987 ( .I0(regs[858]), .I1(wdata[26]), .S(n1217), .Z(n491) );
  CKMUX2V2_8TH40 U988 ( .I0(regs[857]), .I1(wdata[25]), .S(n1217), .Z(n490) );
  CKMUX2V2_8TH40 U989 ( .I0(regs[856]), .I1(wdata[24]), .S(n1217), .Z(n489) );
  CKMUX2V2_8TH40 U990 ( .I0(regs[855]), .I1(wdata[23]), .S(n1217), .Z(n488) );
  CKMUX2V2_8TH40 U991 ( .I0(regs[854]), .I1(wdata[22]), .S(n1217), .Z(n487) );
  CKMUX2V2_8TH40 U992 ( .I0(regs[853]), .I1(wdata[21]), .S(n1217), .Z(n486) );
  CKMUX2V2_8TH40 U993 ( .I0(regs[852]), .I1(wdata[20]), .S(n1217), .Z(n485) );
  CKMUX2V2_8TH40 U994 ( .I0(regs[851]), .I1(wdata[19]), .S(n1217), .Z(n484) );
  CKMUX2V2_8TH40 U995 ( .I0(regs[850]), .I1(wdata[18]), .S(n1217), .Z(n483) );
  CKMUX2V2_8TH40 U996 ( .I0(regs[849]), .I1(wdata[17]), .S(n1217), .Z(n482) );
  CKMUX2V2_8TH40 U997 ( .I0(regs[848]), .I1(wdata[16]), .S(n1217), .Z(n481) );
  CKMUX2V2_8TH40 U998 ( .I0(regs[847]), .I1(wdata[15]), .S(n1217), .Z(n480) );
  CKMUX2V2_8TH40 U999 ( .I0(regs[846]), .I1(wdata[14]), .S(n1217), .Z(n479) );
  CKMUX2V2_8TH40 U1000 ( .I0(regs[845]), .I1(wdata[13]), .S(n1217), .Z(n478)
         );
  CKMUX2V2_8TH40 U1001 ( .I0(regs[844]), .I1(wdata[12]), .S(n1217), .Z(n477)
         );
  CKMUX2V2_8TH40 U1002 ( .I0(regs[843]), .I1(wdata[11]), .S(n1217), .Z(n476)
         );
  CKMUX2V2_8TH40 U1003 ( .I0(regs[842]), .I1(wdata[10]), .S(n1217), .Z(n475)
         );
  CKMUX2V2_8TH40 U1004 ( .I0(regs[841]), .I1(wdata[9]), .S(n1217), .Z(n474) );
  CKMUX2V2_8TH40 U1005 ( .I0(regs[840]), .I1(wdata[8]), .S(n1217), .Z(n473) );
  CKMUX2V2_8TH40 U1006 ( .I0(regs[839]), .I1(wdata[7]), .S(n1217), .Z(n472) );
  CKMUX2V2_8TH40 U1007 ( .I0(regs[838]), .I1(wdata[6]), .S(n1217), .Z(n471) );
  CKMUX2V2_8TH40 U1008 ( .I0(regs[837]), .I1(wdata[5]), .S(n1217), .Z(n470) );
  CKMUX2V2_8TH40 U1009 ( .I0(regs[836]), .I1(wdata[4]), .S(n1217), .Z(n469) );
  CKMUX2V2_8TH40 U1010 ( .I0(regs[835]), .I1(wdata[3]), .S(n1217), .Z(n468) );
  CKMUX2V2_8TH40 U1011 ( .I0(regs[834]), .I1(wdata[2]), .S(n1217), .Z(n467) );
  CKMUX2V2_8TH40 U1012 ( .I0(regs[833]), .I1(wdata[1]), .S(n1217), .Z(n466) );
  CKMUX2V2_8TH40 U1013 ( .I0(regs[832]), .I1(wdata[0]), .S(n1217), .Z(n465) );
  CKMUX2V2_8TH40 U1014 ( .I0(regs[831]), .I1(wdata[31]), .S(n1218), .Z(n464)
         );
  CKMUX2V2_8TH40 U1015 ( .I0(regs[830]), .I1(wdata[30]), .S(n1218), .Z(n463)
         );
  CKMUX2V2_8TH40 U1016 ( .I0(regs[829]), .I1(wdata[29]), .S(n1218), .Z(n462)
         );
  CKMUX2V2_8TH40 U1017 ( .I0(regs[828]), .I1(wdata[28]), .S(n1218), .Z(n461)
         );
  CKMUX2V2_8TH40 U1018 ( .I0(regs[827]), .I1(wdata[27]), .S(n1218), .Z(n460)
         );
  CKMUX2V2_8TH40 U1019 ( .I0(regs[826]), .I1(wdata[26]), .S(n1218), .Z(n459)
         );
  CKMUX2V2_8TH40 U1020 ( .I0(regs[825]), .I1(wdata[25]), .S(n1218), .Z(n458)
         );
  CKMUX2V2_8TH40 U1021 ( .I0(regs[824]), .I1(wdata[24]), .S(n1218), .Z(n457)
         );
  CKMUX2V2_8TH40 U1022 ( .I0(regs[823]), .I1(wdata[23]), .S(n1218), .Z(n456)
         );
  CKMUX2V2_8TH40 U1023 ( .I0(regs[822]), .I1(wdata[22]), .S(n1218), .Z(n455)
         );
  CKMUX2V2_8TH40 U1024 ( .I0(regs[821]), .I1(wdata[21]), .S(n1218), .Z(n454)
         );
  CKMUX2V2_8TH40 U1025 ( .I0(regs[820]), .I1(wdata[20]), .S(n1218), .Z(n453)
         );
  CKMUX2V2_8TH40 U1026 ( .I0(regs[819]), .I1(wdata[19]), .S(n1218), .Z(n452)
         );
  CKMUX2V2_8TH40 U1027 ( .I0(regs[818]), .I1(wdata[18]), .S(n1218), .Z(n451)
         );
  CKMUX2V2_8TH40 U1028 ( .I0(regs[817]), .I1(wdata[17]), .S(n1218), .Z(n450)
         );
  CKMUX2V2_8TH40 U1029 ( .I0(regs[816]), .I1(wdata[16]), .S(n1218), .Z(n449)
         );
  CKMUX2V2_8TH40 U1030 ( .I0(regs[815]), .I1(wdata[15]), .S(n1218), .Z(n448)
         );
  CKMUX2V2_8TH40 U1031 ( .I0(regs[814]), .I1(wdata[14]), .S(n1218), .Z(n447)
         );
  CKMUX2V2_8TH40 U1032 ( .I0(regs[813]), .I1(wdata[13]), .S(n1218), .Z(n446)
         );
  CKMUX2V2_8TH40 U1033 ( .I0(regs[812]), .I1(wdata[12]), .S(n1218), .Z(n445)
         );
  CKMUX2V2_8TH40 U1034 ( .I0(regs[811]), .I1(wdata[11]), .S(n1218), .Z(n444)
         );
  CKMUX2V2_8TH40 U1035 ( .I0(regs[810]), .I1(wdata[10]), .S(n1218), .Z(n443)
         );
  CKMUX2V2_8TH40 U1036 ( .I0(regs[809]), .I1(wdata[9]), .S(n1218), .Z(n442) );
  CKMUX2V2_8TH40 U1037 ( .I0(regs[808]), .I1(wdata[8]), .S(n1218), .Z(n441) );
  CKMUX2V2_8TH40 U1038 ( .I0(regs[807]), .I1(wdata[7]), .S(n1218), .Z(n440) );
  CKMUX2V2_8TH40 U1039 ( .I0(regs[806]), .I1(wdata[6]), .S(n1218), .Z(n439) );
  CKMUX2V2_8TH40 U1040 ( .I0(regs[805]), .I1(wdata[5]), .S(n1218), .Z(n438) );
  CKMUX2V2_8TH40 U1041 ( .I0(regs[804]), .I1(wdata[4]), .S(n1218), .Z(n437) );
  CKMUX2V2_8TH40 U1042 ( .I0(regs[803]), .I1(wdata[3]), .S(n1218), .Z(n436) );
  CKMUX2V2_8TH40 U1043 ( .I0(regs[802]), .I1(wdata[2]), .S(n1218), .Z(n435) );
  CKMUX2V2_8TH40 U1044 ( .I0(regs[801]), .I1(wdata[1]), .S(n1218), .Z(n434) );
  CKMUX2V2_8TH40 U1045 ( .I0(regs[800]), .I1(wdata[0]), .S(n1218), .Z(n433) );
  CKMUX2V2_8TH40 U1046 ( .I0(regs[799]), .I1(wdata[31]), .S(n1219), .Z(n432)
         );
  CKMUX2V2_8TH40 U1047 ( .I0(regs[798]), .I1(wdata[30]), .S(n1219), .Z(n431)
         );
  CKMUX2V2_8TH40 U1048 ( .I0(regs[797]), .I1(wdata[29]), .S(n1219), .Z(n430)
         );
  CKMUX2V2_8TH40 U1049 ( .I0(regs[796]), .I1(wdata[28]), .S(n1219), .Z(n429)
         );
  CKMUX2V2_8TH40 U1050 ( .I0(regs[795]), .I1(wdata[27]), .S(n1219), .Z(n428)
         );
  CKMUX2V2_8TH40 U1051 ( .I0(regs[794]), .I1(wdata[26]), .S(n1219), .Z(n427)
         );
  CKMUX2V2_8TH40 U1052 ( .I0(regs[793]), .I1(wdata[25]), .S(n1219), .Z(n426)
         );
  CKMUX2V2_8TH40 U1053 ( .I0(regs[792]), .I1(wdata[24]), .S(n1219), .Z(n425)
         );
  CKMUX2V2_8TH40 U1054 ( .I0(regs[791]), .I1(wdata[23]), .S(n1219), .Z(n424)
         );
  CKMUX2V2_8TH40 U1055 ( .I0(regs[790]), .I1(wdata[22]), .S(n1219), .Z(n423)
         );
  CKMUX2V2_8TH40 U1056 ( .I0(regs[789]), .I1(wdata[21]), .S(n1219), .Z(n422)
         );
  CKMUX2V2_8TH40 U1057 ( .I0(regs[788]), .I1(wdata[20]), .S(n1219), .Z(n421)
         );
  CKMUX2V2_8TH40 U1058 ( .I0(regs[787]), .I1(wdata[19]), .S(n1219), .Z(n420)
         );
  CKMUX2V2_8TH40 U1059 ( .I0(regs[786]), .I1(wdata[18]), .S(n1219), .Z(n419)
         );
  CKMUX2V2_8TH40 U1060 ( .I0(regs[785]), .I1(wdata[17]), .S(n1219), .Z(n418)
         );
  CKMUX2V2_8TH40 U1061 ( .I0(regs[784]), .I1(wdata[16]), .S(n1219), .Z(n417)
         );
  CKMUX2V2_8TH40 U1062 ( .I0(regs[783]), .I1(wdata[15]), .S(n1219), .Z(n416)
         );
  CKMUX2V2_8TH40 U1063 ( .I0(regs[782]), .I1(wdata[14]), .S(n1219), .Z(n415)
         );
  CKMUX2V2_8TH40 U1064 ( .I0(regs[781]), .I1(wdata[13]), .S(n1219), .Z(n414)
         );
  CKMUX2V2_8TH40 U1065 ( .I0(regs[780]), .I1(wdata[12]), .S(n1219), .Z(n413)
         );
  CKMUX2V2_8TH40 U1066 ( .I0(regs[779]), .I1(wdata[11]), .S(n1219), .Z(n412)
         );
  CKMUX2V2_8TH40 U1067 ( .I0(regs[778]), .I1(wdata[10]), .S(n1219), .Z(n411)
         );
  CKMUX2V2_8TH40 U1068 ( .I0(regs[777]), .I1(wdata[9]), .S(n1219), .Z(n410) );
  CKMUX2V2_8TH40 U1069 ( .I0(regs[776]), .I1(wdata[8]), .S(n1219), .Z(n409) );
  CKMUX2V2_8TH40 U1070 ( .I0(regs[775]), .I1(wdata[7]), .S(n1219), .Z(n408) );
  CKMUX2V2_8TH40 U1071 ( .I0(regs[774]), .I1(wdata[6]), .S(n1219), .Z(n407) );
  CKMUX2V2_8TH40 U1072 ( .I0(regs[773]), .I1(wdata[5]), .S(n1219), .Z(n406) );
  CKMUX2V2_8TH40 U1073 ( .I0(regs[772]), .I1(wdata[4]), .S(n1219), .Z(n405) );
  CKMUX2V2_8TH40 U1074 ( .I0(regs[771]), .I1(wdata[3]), .S(n1219), .Z(n404) );
  CKMUX2V2_8TH40 U1075 ( .I0(regs[770]), .I1(wdata[2]), .S(n1219), .Z(n403) );
  CKMUX2V2_8TH40 U1076 ( .I0(regs[769]), .I1(wdata[1]), .S(n1219), .Z(n402) );
  CKMUX2V2_8TH40 U1077 ( .I0(regs[768]), .I1(wdata[0]), .S(n1219), .Z(n401) );
  NAND3V0P5_8TH40 U1078 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1205) );
  CKMUX2V2_8TH40 U1079 ( .I0(regs[671]), .I1(wdata[31]), .S(n1224), .Z(n400)
         );
  CKMUX2V2_8TH40 U1080 ( .I0(regs[670]), .I1(wdata[30]), .S(n1224), .Z(n399)
         );
  CKMUX2V2_8TH40 U1081 ( .I0(regs[669]), .I1(wdata[29]), .S(n1224), .Z(n398)
         );
  CKMUX2V2_8TH40 U1082 ( .I0(regs[668]), .I1(wdata[28]), .S(n1224), .Z(n397)
         );
  CKMUX2V2_8TH40 U1083 ( .I0(regs[667]), .I1(wdata[27]), .S(n1224), .Z(n396)
         );
  CKMUX2V2_8TH40 U1084 ( .I0(regs[666]), .I1(wdata[26]), .S(n1224), .Z(n395)
         );
  CKMUX2V2_8TH40 U1085 ( .I0(regs[665]), .I1(wdata[25]), .S(n1224), .Z(n394)
         );
  CKMUX2V2_8TH40 U1086 ( .I0(regs[664]), .I1(wdata[24]), .S(n1224), .Z(n393)
         );
  CKMUX2V2_8TH40 U1087 ( .I0(regs[663]), .I1(wdata[23]), .S(n1224), .Z(n392)
         );
  CKMUX2V2_8TH40 U1088 ( .I0(regs[662]), .I1(wdata[22]), .S(n1224), .Z(n391)
         );
  CKMUX2V2_8TH40 U1089 ( .I0(regs[661]), .I1(wdata[21]), .S(n1224), .Z(n390)
         );
  CKMUX2V2_8TH40 U1090 ( .I0(regs[660]), .I1(wdata[20]), .S(n1224), .Z(n389)
         );
  CKMUX2V2_8TH40 U1091 ( .I0(regs[659]), .I1(wdata[19]), .S(n1224), .Z(n388)
         );
  CKMUX2V2_8TH40 U1092 ( .I0(regs[658]), .I1(wdata[18]), .S(n1224), .Z(n387)
         );
  CKMUX2V2_8TH40 U1093 ( .I0(regs[657]), .I1(wdata[17]), .S(n1224), .Z(n386)
         );
  CKMUX2V2_8TH40 U1094 ( .I0(regs[656]), .I1(wdata[16]), .S(n1224), .Z(n385)
         );
  CKMUX2V2_8TH40 U1095 ( .I0(regs[655]), .I1(wdata[15]), .S(n1224), .Z(n384)
         );
  CKMUX2V2_8TH40 U1096 ( .I0(regs[654]), .I1(wdata[14]), .S(n1224), .Z(n383)
         );
  CKMUX2V2_8TH40 U1097 ( .I0(regs[653]), .I1(wdata[13]), .S(n1224), .Z(n382)
         );
  CKMUX2V2_8TH40 U1098 ( .I0(regs[652]), .I1(wdata[12]), .S(n1224), .Z(n381)
         );
  CKMUX2V2_8TH40 U1099 ( .I0(regs[651]), .I1(wdata[11]), .S(n1224), .Z(n380)
         );
  CKMUX2V2_8TH40 U1100 ( .I0(regs[650]), .I1(wdata[10]), .S(n1224), .Z(n379)
         );
  CKMUX2V2_8TH40 U1101 ( .I0(regs[649]), .I1(wdata[9]), .S(n1224), .Z(n378) );
  CKMUX2V2_8TH40 U1102 ( .I0(regs[648]), .I1(wdata[8]), .S(n1224), .Z(n377) );
  CKMUX2V2_8TH40 U1103 ( .I0(regs[647]), .I1(wdata[7]), .S(n1224), .Z(n376) );
  CKMUX2V2_8TH40 U1104 ( .I0(regs[646]), .I1(wdata[6]), .S(n1224), .Z(n375) );
  CKMUX2V2_8TH40 U1105 ( .I0(regs[645]), .I1(wdata[5]), .S(n1224), .Z(n374) );
  CKMUX2V2_8TH40 U1106 ( .I0(regs[644]), .I1(wdata[4]), .S(n1224), .Z(n373) );
  CKMUX2V2_8TH40 U1107 ( .I0(regs[643]), .I1(wdata[3]), .S(n1224), .Z(n372) );
  CKMUX2V2_8TH40 U1108 ( .I0(regs[642]), .I1(wdata[2]), .S(n1224), .Z(n371) );
  CKMUX2V2_8TH40 U1109 ( .I0(regs[641]), .I1(wdata[1]), .S(n1224), .Z(n370) );
  CKMUX2V2_8TH40 U1110 ( .I0(regs[640]), .I1(wdata[0]), .S(n1224), .Z(n369) );
  CKMUX2V2_8TH40 U1111 ( .I0(regs[607]), .I1(wdata[31]), .S(n1225), .Z(n368)
         );
  CKMUX2V2_8TH40 U1112 ( .I0(regs[606]), .I1(wdata[30]), .S(n1225), .Z(n367)
         );
  CKMUX2V2_8TH40 U1113 ( .I0(regs[605]), .I1(wdata[29]), .S(n1225), .Z(n366)
         );
  CKMUX2V2_8TH40 U1114 ( .I0(regs[604]), .I1(wdata[28]), .S(n1225), .Z(n365)
         );
  CKMUX2V2_8TH40 U1115 ( .I0(regs[603]), .I1(wdata[27]), .S(n1225), .Z(n364)
         );
  CKMUX2V2_8TH40 U1116 ( .I0(regs[602]), .I1(wdata[26]), .S(n1225), .Z(n363)
         );
  CKMUX2V2_8TH40 U1117 ( .I0(regs[601]), .I1(wdata[25]), .S(n1225), .Z(n362)
         );
  CKMUX2V2_8TH40 U1118 ( .I0(regs[600]), .I1(wdata[24]), .S(n1225), .Z(n361)
         );
  CKMUX2V2_8TH40 U1119 ( .I0(regs[599]), .I1(wdata[23]), .S(n1225), .Z(n360)
         );
  CKMUX2V2_8TH40 U1120 ( .I0(regs[598]), .I1(wdata[22]), .S(n1225), .Z(n359)
         );
  CKMUX2V2_8TH40 U1121 ( .I0(regs[597]), .I1(wdata[21]), .S(n1225), .Z(n358)
         );
  CKMUX2V2_8TH40 U1122 ( .I0(regs[596]), .I1(wdata[20]), .S(n1225), .Z(n357)
         );
  CKMUX2V2_8TH40 U1123 ( .I0(regs[595]), .I1(wdata[19]), .S(n1225), .Z(n356)
         );
  CKMUX2V2_8TH40 U1124 ( .I0(regs[594]), .I1(wdata[18]), .S(n1225), .Z(n355)
         );
  CKMUX2V2_8TH40 U1125 ( .I0(regs[593]), .I1(wdata[17]), .S(n1225), .Z(n354)
         );
  CKMUX2V2_8TH40 U1126 ( .I0(regs[592]), .I1(wdata[16]), .S(n1225), .Z(n353)
         );
  CKMUX2V2_8TH40 U1127 ( .I0(regs[591]), .I1(wdata[15]), .S(n1225), .Z(n352)
         );
  CKMUX2V2_8TH40 U1128 ( .I0(regs[590]), .I1(wdata[14]), .S(n1225), .Z(n351)
         );
  CKMUX2V2_8TH40 U1129 ( .I0(regs[589]), .I1(wdata[13]), .S(n1225), .Z(n350)
         );
  CKMUX2V2_8TH40 U1130 ( .I0(regs[588]), .I1(wdata[12]), .S(n1225), .Z(n349)
         );
  CKMUX2V2_8TH40 U1131 ( .I0(regs[587]), .I1(wdata[11]), .S(n1225), .Z(n348)
         );
  CKMUX2V2_8TH40 U1132 ( .I0(regs[586]), .I1(wdata[10]), .S(n1225), .Z(n347)
         );
  CKMUX2V2_8TH40 U1133 ( .I0(regs[585]), .I1(wdata[9]), .S(n1225), .Z(n346) );
  CKMUX2V2_8TH40 U1134 ( .I0(regs[584]), .I1(wdata[8]), .S(n1225), .Z(n345) );
  CKMUX2V2_8TH40 U1135 ( .I0(regs[583]), .I1(wdata[7]), .S(n1225), .Z(n344) );
  CKMUX2V2_8TH40 U1136 ( .I0(regs[582]), .I1(wdata[6]), .S(n1225), .Z(n343) );
  CKMUX2V2_8TH40 U1137 ( .I0(regs[581]), .I1(wdata[5]), .S(n1225), .Z(n342) );
  CKMUX2V2_8TH40 U1138 ( .I0(regs[580]), .I1(wdata[4]), .S(n1225), .Z(n341) );
  CKMUX2V2_8TH40 U1139 ( .I0(regs[579]), .I1(wdata[3]), .S(n1225), .Z(n340) );
  CKMUX2V2_8TH40 U1140 ( .I0(regs[578]), .I1(wdata[2]), .S(n1225), .Z(n339) );
  CKMUX2V2_8TH40 U1141 ( .I0(regs[577]), .I1(wdata[1]), .S(n1225), .Z(n338) );
  CKMUX2V2_8TH40 U1142 ( .I0(regs[576]), .I1(wdata[0]), .S(n1225), .Z(n337) );
  CKMUX2V2_8TH40 U1143 ( .I0(regs[575]), .I1(wdata[31]), .S(n1226), .Z(n336)
         );
  CKMUX2V2_8TH40 U1144 ( .I0(regs[574]), .I1(wdata[30]), .S(n1226), .Z(n335)
         );
  CKMUX2V2_8TH40 U1145 ( .I0(regs[573]), .I1(wdata[29]), .S(n1226), .Z(n334)
         );
  CKMUX2V2_8TH40 U1146 ( .I0(regs[572]), .I1(wdata[28]), .S(n1226), .Z(n333)
         );
  CKMUX2V2_8TH40 U1147 ( .I0(regs[571]), .I1(wdata[27]), .S(n1226), .Z(n332)
         );
  CKMUX2V2_8TH40 U1148 ( .I0(regs[570]), .I1(wdata[26]), .S(n1226), .Z(n331)
         );
  CKMUX2V2_8TH40 U1149 ( .I0(regs[569]), .I1(wdata[25]), .S(n1226), .Z(n330)
         );
  CKMUX2V2_8TH40 U1150 ( .I0(regs[568]), .I1(wdata[24]), .S(n1226), .Z(n329)
         );
  CKMUX2V2_8TH40 U1151 ( .I0(regs[567]), .I1(wdata[23]), .S(n1226), .Z(n328)
         );
  CKMUX2V2_8TH40 U1152 ( .I0(regs[566]), .I1(wdata[22]), .S(n1226), .Z(n327)
         );
  CKMUX2V2_8TH40 U1153 ( .I0(regs[565]), .I1(wdata[21]), .S(n1226), .Z(n326)
         );
  CKMUX2V2_8TH40 U1154 ( .I0(regs[564]), .I1(wdata[20]), .S(n1226), .Z(n325)
         );
  CKMUX2V2_8TH40 U1155 ( .I0(regs[563]), .I1(wdata[19]), .S(n1226), .Z(n324)
         );
  CKMUX2V2_8TH40 U1156 ( .I0(regs[562]), .I1(wdata[18]), .S(n1226), .Z(n323)
         );
  CKMUX2V2_8TH40 U1157 ( .I0(regs[561]), .I1(wdata[17]), .S(n1226), .Z(n322)
         );
  CKMUX2V2_8TH40 U1158 ( .I0(regs[560]), .I1(wdata[16]), .S(n1226), .Z(n321)
         );
  CKMUX2V2_8TH40 U1159 ( .I0(regs[559]), .I1(wdata[15]), .S(n1226), .Z(n320)
         );
  CKMUX2V2_8TH40 U1160 ( .I0(regs[558]), .I1(wdata[14]), .S(n1226), .Z(n319)
         );
  CKMUX2V2_8TH40 U1161 ( .I0(regs[557]), .I1(wdata[13]), .S(n1226), .Z(n318)
         );
  CKMUX2V2_8TH40 U1162 ( .I0(regs[556]), .I1(wdata[12]), .S(n1226), .Z(n317)
         );
  CKMUX2V2_8TH40 U1163 ( .I0(regs[555]), .I1(wdata[11]), .S(n1226), .Z(n316)
         );
  CKMUX2V2_8TH40 U1164 ( .I0(regs[554]), .I1(wdata[10]), .S(n1226), .Z(n315)
         );
  CKMUX2V2_8TH40 U1165 ( .I0(regs[553]), .I1(wdata[9]), .S(n1226), .Z(n314) );
  CKMUX2V2_8TH40 U1166 ( .I0(regs[552]), .I1(wdata[8]), .S(n1226), .Z(n313) );
  CKMUX2V2_8TH40 U1167 ( .I0(regs[551]), .I1(wdata[7]), .S(n1226), .Z(n312) );
  CKMUX2V2_8TH40 U1168 ( .I0(regs[550]), .I1(wdata[6]), .S(n1226), .Z(n311) );
  CKMUX2V2_8TH40 U1169 ( .I0(regs[549]), .I1(wdata[5]), .S(n1226), .Z(n310) );
  CKMUX2V2_8TH40 U1170 ( .I0(regs[548]), .I1(wdata[4]), .S(n1226), .Z(n309) );
  CKMUX2V2_8TH40 U1171 ( .I0(regs[547]), .I1(wdata[3]), .S(n1226), .Z(n308) );
  CKMUX2V2_8TH40 U1172 ( .I0(regs[546]), .I1(wdata[2]), .S(n1226), .Z(n307) );
  CKMUX2V2_8TH40 U1173 ( .I0(regs[545]), .I1(wdata[1]), .S(n1226), .Z(n306) );
  CKMUX2V2_8TH40 U1174 ( .I0(regs[544]), .I1(wdata[0]), .S(n1226), .Z(n305) );
  CKMUX2V2_8TH40 U1175 ( .I0(regs[543]), .I1(wdata[31]), .S(n1227), .Z(n304)
         );
  CKMUX2V2_8TH40 U1176 ( .I0(regs[542]), .I1(wdata[30]), .S(n1227), .Z(n303)
         );
  CKMUX2V2_8TH40 U1177 ( .I0(regs[541]), .I1(wdata[29]), .S(n1227), .Z(n302)
         );
  CKMUX2V2_8TH40 U1178 ( .I0(regs[540]), .I1(wdata[28]), .S(n1227), .Z(n301)
         );
  CKMUX2V2_8TH40 U1179 ( .I0(regs[539]), .I1(wdata[27]), .S(n1227), .Z(n300)
         );
  CKMUX2V2_8TH40 U1180 ( .I0(regs[538]), .I1(wdata[26]), .S(n1227), .Z(n299)
         );
  CKMUX2V2_8TH40 U1181 ( .I0(regs[537]), .I1(wdata[25]), .S(n1227), .Z(n298)
         );
  CKMUX2V2_8TH40 U1182 ( .I0(regs[536]), .I1(wdata[24]), .S(n1227), .Z(n297)
         );
  CKMUX2V2_8TH40 U1183 ( .I0(regs[535]), .I1(wdata[23]), .S(n1227), .Z(n296)
         );
  CKMUX2V2_8TH40 U1184 ( .I0(regs[534]), .I1(wdata[22]), .S(n1227), .Z(n295)
         );
  CKMUX2V2_8TH40 U1185 ( .I0(regs[533]), .I1(wdata[21]), .S(n1227), .Z(n294)
         );
  CKMUX2V2_8TH40 U1186 ( .I0(regs[532]), .I1(wdata[20]), .S(n1227), .Z(n293)
         );
  CKMUX2V2_8TH40 U1187 ( .I0(regs[531]), .I1(wdata[19]), .S(n1227), .Z(n292)
         );
  CKMUX2V2_8TH40 U1188 ( .I0(regs[530]), .I1(wdata[18]), .S(n1227), .Z(n291)
         );
  CKMUX2V2_8TH40 U1189 ( .I0(regs[529]), .I1(wdata[17]), .S(n1227), .Z(n290)
         );
  CKMUX2V2_8TH40 U1190 ( .I0(regs[528]), .I1(wdata[16]), .S(n1227), .Z(n289)
         );
  CKMUX2V2_8TH40 U1191 ( .I0(regs[527]), .I1(wdata[15]), .S(n1227), .Z(n288)
         );
  CKMUX2V2_8TH40 U1192 ( .I0(regs[526]), .I1(wdata[14]), .S(n1227), .Z(n287)
         );
  CKMUX2V2_8TH40 U1193 ( .I0(regs[525]), .I1(wdata[13]), .S(n1227), .Z(n286)
         );
  CKMUX2V2_8TH40 U1194 ( .I0(regs[524]), .I1(wdata[12]), .S(n1227), .Z(n285)
         );
  CKMUX2V2_8TH40 U1195 ( .I0(regs[523]), .I1(wdata[11]), .S(n1227), .Z(n284)
         );
  CKMUX2V2_8TH40 U1196 ( .I0(regs[522]), .I1(wdata[10]), .S(n1227), .Z(n283)
         );
  CKMUX2V2_8TH40 U1197 ( .I0(regs[521]), .I1(wdata[9]), .S(n1227), .Z(n282) );
  CKMUX2V2_8TH40 U1198 ( .I0(regs[520]), .I1(wdata[8]), .S(n1227), .Z(n281) );
  CKMUX2V2_8TH40 U1199 ( .I0(regs[519]), .I1(wdata[7]), .S(n1227), .Z(n280) );
  CKMUX2V2_8TH40 U1200 ( .I0(regs[518]), .I1(wdata[6]), .S(n1227), .Z(n279) );
  CKMUX2V2_8TH40 U1201 ( .I0(regs[517]), .I1(wdata[5]), .S(n1227), .Z(n278) );
  CKMUX2V2_8TH40 U1202 ( .I0(regs[516]), .I1(wdata[4]), .S(n1227), .Z(n277) );
  CKMUX2V2_8TH40 U1203 ( .I0(regs[515]), .I1(wdata[3]), .S(n1227), .Z(n276) );
  CKMUX2V2_8TH40 U1204 ( .I0(regs[514]), .I1(wdata[2]), .S(n1227), .Z(n275) );
  CKMUX2V2_8TH40 U1205 ( .I0(regs[513]), .I1(wdata[1]), .S(n1227), .Z(n274) );
  CKMUX2V2_8TH40 U1206 ( .I0(regs[512]), .I1(wdata[0]), .S(n1227), .Z(n273) );
  NAND3V0P5_8TH40 U1207 ( .A1(waddr[3]), .A2(n1222), .A3(n1223), .ZN(n1208) );
  CLKNV1_8TH40 U1208 ( .I(waddr[4]), .ZN(n1222) );
  CKMUX2V2_8TH40 U1209 ( .I0(regs[287]), .I1(wdata[31]), .S(n1228), .Z(n272)
         );
  CKMUX2V2_8TH40 U1210 ( .I0(regs[286]), .I1(wdata[30]), .S(n1228), .Z(n271)
         );
  CKMUX2V2_8TH40 U1211 ( .I0(regs[285]), .I1(wdata[29]), .S(n1228), .Z(n270)
         );
  CKMUX2V2_8TH40 U1212 ( .I0(regs[284]), .I1(wdata[28]), .S(n1228), .Z(n269)
         );
  CKMUX2V2_8TH40 U1213 ( .I0(regs[283]), .I1(wdata[27]), .S(n1228), .Z(n268)
         );
  CKMUX2V2_8TH40 U1214 ( .I0(regs[282]), .I1(wdata[26]), .S(n1228), .Z(n267)
         );
  CKMUX2V2_8TH40 U1215 ( .I0(regs[281]), .I1(wdata[25]), .S(n1228), .Z(n266)
         );
  CKMUX2V2_8TH40 U1216 ( .I0(regs[280]), .I1(wdata[24]), .S(n1228), .Z(n265)
         );
  CKMUX2V2_8TH40 U1217 ( .I0(regs[279]), .I1(wdata[23]), .S(n1228), .Z(n264)
         );
  CKMUX2V2_8TH40 U1218 ( .I0(regs[278]), .I1(wdata[22]), .S(n1228), .Z(n263)
         );
  CKMUX2V2_8TH40 U1219 ( .I0(regs[277]), .I1(wdata[21]), .S(n1228), .Z(n262)
         );
  CKMUX2V2_8TH40 U1220 ( .I0(regs[276]), .I1(wdata[20]), .S(n1228), .Z(n261)
         );
  CKMUX2V2_8TH40 U1221 ( .I0(regs[275]), .I1(wdata[19]), .S(n1228), .Z(n260)
         );
  CKMUX2V2_8TH40 U1222 ( .I0(regs[274]), .I1(wdata[18]), .S(n1228), .Z(n259)
         );
  CKMUX2V2_8TH40 U1223 ( .I0(regs[273]), .I1(wdata[17]), .S(n1228), .Z(n258)
         );
  CKMUX2V2_8TH40 U1224 ( .I0(regs[272]), .I1(wdata[16]), .S(n1228), .Z(n257)
         );
  CKMUX2V2_8TH40 U1225 ( .I0(regs[271]), .I1(wdata[15]), .S(n1228), .Z(n256)
         );
  CKMUX2V2_8TH40 U1226 ( .I0(regs[270]), .I1(wdata[14]), .S(n1228), .Z(n255)
         );
  CKMUX2V2_8TH40 U1227 ( .I0(regs[269]), .I1(wdata[13]), .S(n1228), .Z(n254)
         );
  CKMUX2V2_8TH40 U1228 ( .I0(regs[268]), .I1(wdata[12]), .S(n1228), .Z(n253)
         );
  CKMUX2V2_8TH40 U1229 ( .I0(regs[267]), .I1(wdata[11]), .S(n1228), .Z(n252)
         );
  CKMUX2V2_8TH40 U1230 ( .I0(regs[266]), .I1(wdata[10]), .S(n1228), .Z(n251)
         );
  CKMUX2V2_8TH40 U1231 ( .I0(regs[265]), .I1(wdata[9]), .S(n1228), .Z(n250) );
  CKMUX2V2_8TH40 U1232 ( .I0(regs[264]), .I1(wdata[8]), .S(n1228), .Z(n249) );
  CKMUX2V2_8TH40 U1233 ( .I0(regs[263]), .I1(wdata[7]), .S(n1228), .Z(n248) );
  CKMUX2V2_8TH40 U1234 ( .I0(regs[262]), .I1(wdata[6]), .S(n1228), .Z(n247) );
  CKMUX2V2_8TH40 U1235 ( .I0(regs[261]), .I1(wdata[5]), .S(n1228), .Z(n246) );
  CKMUX2V2_8TH40 U1236 ( .I0(regs[260]), .I1(wdata[4]), .S(n1228), .Z(n245) );
  CKMUX2V2_8TH40 U1237 ( .I0(regs[259]), .I1(wdata[3]), .S(n1228), .Z(n244) );
  CKMUX2V2_8TH40 U1238 ( .I0(regs[258]), .I1(wdata[2]), .S(n1228), .Z(n243) );
  CKMUX2V2_8TH40 U1239 ( .I0(regs[257]), .I1(wdata[1]), .S(n1228), .Z(n242) );
  CKMUX2V2_8TH40 U1240 ( .I0(regs[256]), .I1(wdata[0]), .S(n1228), .Z(n241) );
  NAND3V0P5_8TH40 U1241 ( .A1(waddr[4]), .A2(n1221), .A3(n1223), .ZN(n1210) );
  CLKNV1_8TH40 U1242 ( .I(waddr[3]), .ZN(n1221) );
  CKMUX2V2_8TH40 U1243 ( .I0(regs[159]), .I1(wdata[31]), .S(n1229), .Z(n240)
         );
  CKMUX2V2_8TH40 U1244 ( .I0(regs[158]), .I1(wdata[30]), .S(n1229), .Z(n239)
         );
  CKMUX2V2_8TH40 U1245 ( .I0(regs[157]), .I1(wdata[29]), .S(n1229), .Z(n238)
         );
  CKMUX2V2_8TH40 U1246 ( .I0(regs[156]), .I1(wdata[28]), .S(n1229), .Z(n237)
         );
  CKMUX2V2_8TH40 U1247 ( .I0(regs[155]), .I1(wdata[27]), .S(n1229), .Z(n236)
         );
  CKMUX2V2_8TH40 U1248 ( .I0(regs[154]), .I1(wdata[26]), .S(n1229), .Z(n235)
         );
  CKMUX2V2_8TH40 U1249 ( .I0(regs[153]), .I1(wdata[25]), .S(n1229), .Z(n234)
         );
  CKMUX2V2_8TH40 U1250 ( .I0(regs[152]), .I1(wdata[24]), .S(n1229), .Z(n233)
         );
  CKMUX2V2_8TH40 U1251 ( .I0(regs[151]), .I1(wdata[23]), .S(n1229), .Z(n232)
         );
  CKMUX2V2_8TH40 U1252 ( .I0(regs[150]), .I1(wdata[22]), .S(n1229), .Z(n231)
         );
  CKMUX2V2_8TH40 U1253 ( .I0(regs[149]), .I1(wdata[21]), .S(n1229), .Z(n230)
         );
  CKMUX2V2_8TH40 U1254 ( .I0(regs[148]), .I1(wdata[20]), .S(n1229), .Z(n229)
         );
  CKMUX2V2_8TH40 U1255 ( .I0(regs[147]), .I1(wdata[19]), .S(n1229), .Z(n228)
         );
  CKMUX2V2_8TH40 U1256 ( .I0(regs[146]), .I1(wdata[18]), .S(n1229), .Z(n227)
         );
  CKMUX2V2_8TH40 U1257 ( .I0(regs[145]), .I1(wdata[17]), .S(n1229), .Z(n226)
         );
  CKMUX2V2_8TH40 U1258 ( .I0(regs[144]), .I1(wdata[16]), .S(n1229), .Z(n225)
         );
  CKMUX2V2_8TH40 U1259 ( .I0(regs[143]), .I1(wdata[15]), .S(n1229), .Z(n224)
         );
  CKMUX2V2_8TH40 U1260 ( .I0(regs[142]), .I1(wdata[14]), .S(n1229), .Z(n223)
         );
  CKMUX2V2_8TH40 U1261 ( .I0(regs[141]), .I1(wdata[13]), .S(n1229), .Z(n222)
         );
  CKMUX2V2_8TH40 U1262 ( .I0(regs[140]), .I1(wdata[12]), .S(n1229), .Z(n221)
         );
  CKMUX2V2_8TH40 U1263 ( .I0(regs[139]), .I1(wdata[11]), .S(n1229), .Z(n220)
         );
  CKMUX2V2_8TH40 U1264 ( .I0(regs[138]), .I1(wdata[10]), .S(n1229), .Z(n219)
         );
  CKMUX2V2_8TH40 U1265 ( .I0(regs[137]), .I1(wdata[9]), .S(n1229), .Z(n218) );
  CKMUX2V2_8TH40 U1266 ( .I0(regs[136]), .I1(wdata[8]), .S(n1229), .Z(n217) );
  CKMUX2V2_8TH40 U1267 ( .I0(regs[135]), .I1(wdata[7]), .S(n1229), .Z(n216) );
  CKMUX2V2_8TH40 U1268 ( .I0(regs[134]), .I1(wdata[6]), .S(n1229), .Z(n215) );
  CKMUX2V2_8TH40 U1269 ( .I0(regs[133]), .I1(wdata[5]), .S(n1229), .Z(n214) );
  CKMUX2V2_8TH40 U1270 ( .I0(regs[132]), .I1(wdata[4]), .S(n1229), .Z(n213) );
  CKMUX2V2_8TH40 U1271 ( .I0(regs[131]), .I1(wdata[3]), .S(n1229), .Z(n212) );
  CKMUX2V2_8TH40 U1272 ( .I0(regs[130]), .I1(wdata[2]), .S(n1229), .Z(n211) );
  CKMUX2V2_8TH40 U1273 ( .I0(regs[129]), .I1(wdata[1]), .S(n1229), .Z(n210) );
  CKMUX2V2_8TH40 U1274 ( .I0(regs[128]), .I1(wdata[0]), .S(n1229), .Z(n209) );
  NOR3V0P5_8TH40 U1275 ( .A1(n1192), .A2(waddr[2]), .A3(n1191), .ZN(n1211) );
  CKMUX2V2_8TH40 U1276 ( .I0(regs[95]), .I1(wdata[31]), .S(n1230), .Z(n208) );
  CKMUX2V2_8TH40 U1277 ( .I0(regs[94]), .I1(wdata[30]), .S(n1230), .Z(n207) );
  CKMUX2V2_8TH40 U1278 ( .I0(regs[93]), .I1(wdata[29]), .S(n1230), .Z(n206) );
  CKMUX2V2_8TH40 U1279 ( .I0(regs[92]), .I1(wdata[28]), .S(n1230), .Z(n205) );
  CKMUX2V2_8TH40 U1280 ( .I0(regs[91]), .I1(wdata[27]), .S(n1230), .Z(n204) );
  CKMUX2V2_8TH40 U1281 ( .I0(regs[90]), .I1(wdata[26]), .S(n1230), .Z(n203) );
  CKMUX2V2_8TH40 U1282 ( .I0(regs[89]), .I1(wdata[25]), .S(n1230), .Z(n202) );
  CKMUX2V2_8TH40 U1283 ( .I0(regs[88]), .I1(wdata[24]), .S(n1230), .Z(n201) );
  CKMUX2V2_8TH40 U1284 ( .I0(regs[87]), .I1(wdata[23]), .S(n1230), .Z(n200) );
  CKMUX2V2_8TH40 U1285 ( .I0(regs[86]), .I1(wdata[22]), .S(n1230), .Z(n199) );
  CKMUX2V2_8TH40 U1286 ( .I0(regs[85]), .I1(wdata[21]), .S(n1230), .Z(n198) );
  CKMUX2V2_8TH40 U1287 ( .I0(regs[84]), .I1(wdata[20]), .S(n1230), .Z(n197) );
  CKMUX2V2_8TH40 U1288 ( .I0(regs[83]), .I1(wdata[19]), .S(n1230), .Z(n196) );
  CKMUX2V2_8TH40 U1289 ( .I0(regs[82]), .I1(wdata[18]), .S(n1230), .Z(n195) );
  CKMUX2V2_8TH40 U1290 ( .I0(regs[81]), .I1(wdata[17]), .S(n1230), .Z(n194) );
  CKMUX2V2_8TH40 U1291 ( .I0(regs[80]), .I1(wdata[16]), .S(n1230), .Z(n193) );
  CKMUX2V2_8TH40 U1292 ( .I0(regs[79]), .I1(wdata[15]), .S(n1230), .Z(n192) );
  CKMUX2V2_8TH40 U1293 ( .I0(regs[78]), .I1(wdata[14]), .S(n1230), .Z(n191) );
  CKMUX2V2_8TH40 U1294 ( .I0(regs[77]), .I1(wdata[13]), .S(n1230), .Z(n190) );
  CKMUX2V2_8TH40 U1295 ( .I0(regs[76]), .I1(wdata[12]), .S(n1230), .Z(n189) );
  CKMUX2V2_8TH40 U1296 ( .I0(regs[75]), .I1(wdata[11]), .S(n1230), .Z(n188) );
  CKMUX2V2_8TH40 U1297 ( .I0(regs[74]), .I1(wdata[10]), .S(n1230), .Z(n187) );
  CKMUX2V2_8TH40 U1298 ( .I0(regs[73]), .I1(wdata[9]), .S(n1230), .Z(n186) );
  CKMUX2V2_8TH40 U1299 ( .I0(regs[72]), .I1(wdata[8]), .S(n1230), .Z(n185) );
  CKMUX2V2_8TH40 U1300 ( .I0(regs[71]), .I1(wdata[7]), .S(n1230), .Z(n184) );
  CKMUX2V2_8TH40 U1301 ( .I0(regs[70]), .I1(wdata[6]), .S(n1230), .Z(n183) );
  CKMUX2V2_8TH40 U1302 ( .I0(regs[69]), .I1(wdata[5]), .S(n1230), .Z(n182) );
  CKMUX2V2_8TH40 U1303 ( .I0(regs[68]), .I1(wdata[4]), .S(n1230), .Z(n181) );
  CKMUX2V2_8TH40 U1304 ( .I0(regs[67]), .I1(wdata[3]), .S(n1230), .Z(n180) );
  CKMUX2V2_8TH40 U1305 ( .I0(regs[66]), .I1(wdata[2]), .S(n1230), .Z(n179) );
  CKMUX2V2_8TH40 U1306 ( .I0(regs[65]), .I1(wdata[1]), .S(n1230), .Z(n178) );
  CKMUX2V2_8TH40 U1307 ( .I0(regs[64]), .I1(wdata[0]), .S(n1230), .Z(n177) );
  NOR3V0P5_8TH40 U1308 ( .A1(n1192), .A2(waddr[1]), .A3(n1215), .ZN(n1212) );
  CKMUX2V2_8TH40 U1309 ( .I0(regs[63]), .I1(wdata[31]), .S(n1231), .Z(n176) );
  CKMUX2V2_8TH40 U1310 ( .I0(regs[62]), .I1(wdata[30]), .S(n1231), .Z(n175) );
  CKMUX2V2_8TH40 U1311 ( .I0(regs[61]), .I1(wdata[29]), .S(n1231), .Z(n174) );
  CKMUX2V2_8TH40 U1312 ( .I0(regs[60]), .I1(wdata[28]), .S(n1231), .Z(n173) );
  CKMUX2V2_8TH40 U1313 ( .I0(regs[59]), .I1(wdata[27]), .S(n1231), .Z(n172) );
  CKMUX2V2_8TH40 U1314 ( .I0(regs[58]), .I1(wdata[26]), .S(n1231), .Z(n171) );
  CKMUX2V2_8TH40 U1315 ( .I0(regs[57]), .I1(wdata[25]), .S(n1231), .Z(n170) );
  CKMUX2V2_8TH40 U1316 ( .I0(regs[56]), .I1(wdata[24]), .S(n1231), .Z(n169) );
  CKMUX2V2_8TH40 U1317 ( .I0(regs[55]), .I1(wdata[23]), .S(n1231), .Z(n168) );
  CKMUX2V2_8TH40 U1318 ( .I0(regs[54]), .I1(wdata[22]), .S(n1231), .Z(n167) );
  CKMUX2V2_8TH40 U1319 ( .I0(regs[53]), .I1(wdata[21]), .S(n1231), .Z(n166) );
  CKMUX2V2_8TH40 U1320 ( .I0(regs[52]), .I1(wdata[20]), .S(n1231), .Z(n165) );
  CKMUX2V2_8TH40 U1321 ( .I0(regs[51]), .I1(wdata[19]), .S(n1231), .Z(n164) );
  CKMUX2V2_8TH40 U1322 ( .I0(regs[50]), .I1(wdata[18]), .S(n1231), .Z(n163) );
  CKMUX2V2_8TH40 U1323 ( .I0(regs[49]), .I1(wdata[17]), .S(n1231), .Z(n162) );
  CKMUX2V2_8TH40 U1324 ( .I0(regs[48]), .I1(wdata[16]), .S(n1231), .Z(n161) );
  CKMUX2V2_8TH40 U1325 ( .I0(regs[47]), .I1(wdata[15]), .S(n1231), .Z(n160) );
  CKMUX2V2_8TH40 U1326 ( .I0(regs[46]), .I1(wdata[14]), .S(n1231), .Z(n159) );
  CKMUX2V2_8TH40 U1327 ( .I0(regs[45]), .I1(wdata[13]), .S(n1231), .Z(n158) );
  CKMUX2V2_8TH40 U1328 ( .I0(regs[44]), .I1(wdata[12]), .S(n1231), .Z(n157) );
  CKMUX2V2_8TH40 U1329 ( .I0(regs[43]), .I1(wdata[11]), .S(n1231), .Z(n156) );
  CKMUX2V2_8TH40 U1330 ( .I0(regs[42]), .I1(wdata[10]), .S(n1231), .Z(n155) );
  CKMUX2V2_8TH40 U1331 ( .I0(regs[41]), .I1(wdata[9]), .S(n1231), .Z(n154) );
  CKMUX2V2_8TH40 U1332 ( .I0(regs[40]), .I1(wdata[8]), .S(n1231), .Z(n153) );
  CKMUX2V2_8TH40 U1333 ( .I0(regs[39]), .I1(wdata[7]), .S(n1231), .Z(n152) );
  CKMUX2V2_8TH40 U1334 ( .I0(regs[38]), .I1(wdata[6]), .S(n1231), .Z(n151) );
  CKMUX2V2_8TH40 U1335 ( .I0(regs[37]), .I1(wdata[5]), .S(n1231), .Z(n150) );
  CKMUX2V2_8TH40 U1336 ( .I0(regs[36]), .I1(wdata[4]), .S(n1231), .Z(n149) );
  CKMUX2V2_8TH40 U1337 ( .I0(regs[35]), .I1(wdata[3]), .S(n1231), .Z(n148) );
  CKMUX2V2_8TH40 U1338 ( .I0(regs[34]), .I1(wdata[2]), .S(n1231), .Z(n147) );
  CKMUX2V2_8TH40 U1339 ( .I0(regs[33]), .I1(wdata[1]), .S(n1231), .Z(n146) );
  CKMUX2V2_8TH40 U1340 ( .I0(regs[32]), .I1(wdata[0]), .S(n1231), .Z(n145) );
  NOR3V0P5_8TH40 U1341 ( .A1(n1191), .A2(waddr[0]), .A3(n1215), .ZN(n1213) );
  CKMUX2V2_8TH40 U1342 ( .I0(regs[31]), .I1(wdata[31]), .S(n1232), .Z(n144) );
  CKMUX2V2_8TH40 U1343 ( .I0(regs[30]), .I1(wdata[30]), .S(n1232), .Z(n143) );
  CKMUX2V2_8TH40 U1344 ( .I0(regs[29]), .I1(wdata[29]), .S(n1232), .Z(n142) );
  CKMUX2V2_8TH40 U1345 ( .I0(regs[28]), .I1(wdata[28]), .S(n1232), .Z(n141) );
  CKMUX2V2_8TH40 U1346 ( .I0(regs[27]), .I1(wdata[27]), .S(n1232), .Z(n140) );
  CKMUX2V2_8TH40 U1347 ( .I0(regs[26]), .I1(wdata[26]), .S(n1232), .Z(n139) );
  CKMUX2V2_8TH40 U1348 ( .I0(regs[25]), .I1(wdata[25]), .S(n1232), .Z(n138) );
  CKMUX2V2_8TH40 U1349 ( .I0(regs[24]), .I1(wdata[24]), .S(n1232), .Z(n137) );
  CKMUX2V2_8TH40 U1350 ( .I0(regs[23]), .I1(wdata[23]), .S(n1232), .Z(n136) );
  CKMUX2V2_8TH40 U1351 ( .I0(regs[22]), .I1(wdata[22]), .S(n1232), .Z(n135) );
  CKMUX2V2_8TH40 U1352 ( .I0(regs[21]), .I1(wdata[21]), .S(n1232), .Z(n134) );
  CKMUX2V2_8TH40 U1353 ( .I0(regs[20]), .I1(wdata[20]), .S(n1232), .Z(n133) );
  CKMUX2V2_8TH40 U1354 ( .I0(regs[19]), .I1(wdata[19]), .S(n1232), .Z(n132) );
  CKMUX2V2_8TH40 U1355 ( .I0(regs[18]), .I1(wdata[18]), .S(n1232), .Z(n131) );
  CKMUX2V2_8TH40 U1356 ( .I0(regs[17]), .I1(wdata[17]), .S(n1232), .Z(n130) );
  CKMUX2V2_8TH40 U1357 ( .I0(regs[16]), .I1(wdata[16]), .S(n1232), .Z(n129) );
  CKMUX2V2_8TH40 U1358 ( .I0(regs[15]), .I1(wdata[15]), .S(n1232), .Z(n128) );
  CKMUX2V2_8TH40 U1359 ( .I0(regs[14]), .I1(wdata[14]), .S(n1232), .Z(n127) );
  CKMUX2V2_8TH40 U1360 ( .I0(regs[13]), .I1(wdata[13]), .S(n1232), .Z(n126) );
  CKMUX2V2_8TH40 U1361 ( .I0(regs[12]), .I1(wdata[12]), .S(n1232), .Z(n125) );
  CKMUX2V2_8TH40 U1362 ( .I0(regs[11]), .I1(wdata[11]), .S(n1232), .Z(n124) );
  CKMUX2V2_8TH40 U1363 ( .I0(regs[10]), .I1(wdata[10]), .S(n1232), .Z(n123) );
  CKMUX2V2_8TH40 U1364 ( .I0(regs[9]), .I1(wdata[9]), .S(n1232), .Z(n122) );
  CKMUX2V2_8TH40 U1365 ( .I0(regs[8]), .I1(wdata[8]), .S(n1232), .Z(n121) );
  CKMUX2V2_8TH40 U1366 ( .I0(regs[7]), .I1(wdata[7]), .S(n1232), .Z(n120) );
  CKMUX2V2_8TH40 U1367 ( .I0(regs[6]), .I1(wdata[6]), .S(n1232), .Z(n119) );
  CKMUX2V2_8TH40 U1368 ( .I0(regs[5]), .I1(wdata[5]), .S(n1232), .Z(n118) );
  CKMUX2V2_8TH40 U1369 ( .I0(regs[4]), .I1(wdata[4]), .S(n1232), .Z(n117) );
  CKMUX2V2_8TH40 U1370 ( .I0(regs[3]), .I1(wdata[3]), .S(n1232), .Z(n116) );
  CKMUX2V2_8TH40 U1371 ( .I0(regs[2]), .I1(wdata[2]), .S(n1232), .Z(n115) );
  CKMUX2V2_8TH40 U1372 ( .I0(regs[1]), .I1(wdata[1]), .S(n1232), .Z(n114) );
  CKMUX2V2_8TH40 U1373 ( .I0(regs[0]), .I1(wdata[0]), .S(n1232), .Z(n113) );
  NAND3V0P5_8TH40 U1374 ( .A1(waddr[3]), .A2(waddr[4]), .A3(n1223), .ZN(n1214)
         );
  INOR2V0_8TH40 U1375 ( .A1(we), .B1(rst), .ZN(n1223) );
  NOR3V0P5_8TH40 U1376 ( .A1(n1191), .A2(n1192), .A3(n1215), .ZN(n1220) );
  CLKNV1_8TH40 U1377 ( .I(waddr[2]), .ZN(n1215) );
  CLKNV1_8TH40 U1378 ( .I(waddr[0]), .ZN(n1192) );
  CLKNV1_8TH40 U1379 ( .I(waddr[1]), .ZN(n1191) );
endmodule


module pipe_reg_idex ( clk, rst, stall_ctrl, id_inst_type, id_inst_class, 
        id_gpr1_data, id_gpr2_data, id_target_gpr, id_gpr_we, id_link_addr, 
        id_inst_delayslot, nxtid_inst_delayslot, id_inst, id_except_type, 
        id_cur_inst_addr, ex_inst_type, ex_inst_class, ex_gpr1_data, 
        ex_gpr2_data, ex_target_gpr, ex_gpr_we, ex_link_addr, 
        ex_inst_delayslot, nxt_inst_delayslot, ex_inst, ex_except_type, 
        ex_cur_inst_addr, flush_BAR );
  input [5:0] stall_ctrl;
  input [7:0] id_inst_type;
  input [2:0] id_inst_class;
  input [31:0] id_gpr1_data;
  input [31:0] id_gpr2_data;
  input [4:0] id_target_gpr;
  input [31:0] id_link_addr;
  input [31:0] id_inst;
  input [31:0] id_except_type;
  input [31:0] id_cur_inst_addr;
  output [7:0] ex_inst_type;
  output [2:0] ex_inst_class;
  output [31:0] ex_gpr1_data;
  output [31:0] ex_gpr2_data;
  output [4:0] ex_target_gpr;
  output [31:0] ex_link_addr;
  output [31:0] ex_inst;
  output [31:0] ex_except_type;
  output [31:0] ex_cur_inst_addr;
  input clk, rst, id_gpr_we, id_inst_delayslot, nxtid_inst_delayslot,
         flush_BAR;
  output ex_gpr_we, ex_inst_delayslot, nxt_inst_delayslot;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n159, n160, n163, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n1, n2, n3, n151, n152, n153, n154, n155, n156, n157,
         n158, n161, n162, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180;

  DQV4_8TH40 ex_inst_reg_15_ ( .D(n198), .CK(clk), .Q(ex_inst[15]) );
  DQV4_8TH40 ex_inst_reg_14_ ( .D(n197), .CK(clk), .Q(ex_inst[14]) );
  DQV4_8TH40 ex_inst_reg_13_ ( .D(n196), .CK(clk), .Q(ex_inst[13]) );
  DQV4_8TH40 ex_inst_reg_12_ ( .D(n195), .CK(clk), .Q(ex_inst[12]) );
  DQV4_8TH40 ex_inst_reg_11_ ( .D(n194), .CK(clk), .Q(ex_inst[11]) );
  DQV4_8TH40 ex_inst_reg_10_ ( .D(n193), .CK(clk), .Q(ex_inst[10]) );
  DQV4_8TH40 ex_inst_reg_9_ ( .D(n192), .CK(clk), .Q(ex_inst[9]) );
  DQV4_8TH40 ex_inst_reg_8_ ( .D(n191), .CK(clk), .Q(ex_inst[8]) );
  DQV4_8TH40 ex_inst_reg_7_ ( .D(n190), .CK(clk), .Q(ex_inst[7]) );
  DQV4_8TH40 ex_inst_reg_6_ ( .D(n189), .CK(clk), .Q(ex_inst[6]) );
  DQV4_8TH40 ex_inst_reg_5_ ( .D(n188), .CK(clk), .Q(ex_inst[5]) );
  DQV4_8TH40 ex_inst_reg_4_ ( .D(n187), .CK(clk), .Q(ex_inst[4]) );
  DQV4_8TH40 ex_inst_reg_3_ ( .D(n186), .CK(clk), .Q(ex_inst[3]) );
  DQV4_8TH40 ex_inst_reg_2_ ( .D(n185), .CK(clk), .Q(ex_inst[2]) );
  DQV4_8TH40 ex_inst_reg_1_ ( .D(n184), .CK(clk), .Q(ex_inst[1]) );
  DQV4_8TH40 ex_inst_reg_0_ ( .D(n183), .CK(clk), .Q(ex_inst[0]) );
  DQV4_8TH40 ex_except_type_reg_12_ ( .D(n163), .CK(clk), .Q(
        ex_except_type[12]) );
  DQV4_8TH40 ex_except_type_reg_9_ ( .D(n160), .CK(clk), .Q(ex_except_type[9])
         );
  DQV4_8TH40 ex_except_type_reg_8_ ( .D(n159), .CK(clk), .Q(ex_except_type[8])
         );
  DQV4_8TH40 ex_cur_inst_addr_reg_31_ ( .D(n150), .CK(clk), .Q(
        ex_cur_inst_addr[31]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_30_ ( .D(n149), .CK(clk), .Q(
        ex_cur_inst_addr[30]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_29_ ( .D(n148), .CK(clk), .Q(
        ex_cur_inst_addr[29]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_28_ ( .D(n147), .CK(clk), .Q(
        ex_cur_inst_addr[28]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_27_ ( .D(n146), .CK(clk), .Q(
        ex_cur_inst_addr[27]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_26_ ( .D(n145), .CK(clk), .Q(
        ex_cur_inst_addr[26]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_25_ ( .D(n144), .CK(clk), .Q(
        ex_cur_inst_addr[25]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_24_ ( .D(n143), .CK(clk), .Q(
        ex_cur_inst_addr[24]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_23_ ( .D(n142), .CK(clk), .Q(
        ex_cur_inst_addr[23]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_22_ ( .D(n141), .CK(clk), .Q(
        ex_cur_inst_addr[22]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_21_ ( .D(n140), .CK(clk), .Q(
        ex_cur_inst_addr[21]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_20_ ( .D(n139), .CK(clk), .Q(
        ex_cur_inst_addr[20]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_19_ ( .D(n138), .CK(clk), .Q(
        ex_cur_inst_addr[19]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_18_ ( .D(n137), .CK(clk), .Q(
        ex_cur_inst_addr[18]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_17_ ( .D(n136), .CK(clk), .Q(
        ex_cur_inst_addr[17]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_16_ ( .D(n135), .CK(clk), .Q(
        ex_cur_inst_addr[16]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_15_ ( .D(n134), .CK(clk), .Q(
        ex_cur_inst_addr[15]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_14_ ( .D(n133), .CK(clk), .Q(
        ex_cur_inst_addr[14]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_13_ ( .D(n132), .CK(clk), .Q(
        ex_cur_inst_addr[13]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_12_ ( .D(n131), .CK(clk), .Q(
        ex_cur_inst_addr[12]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_11_ ( .D(n130), .CK(clk), .Q(
        ex_cur_inst_addr[11]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_10_ ( .D(n129), .CK(clk), .Q(
        ex_cur_inst_addr[10]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_9_ ( .D(n128), .CK(clk), .Q(
        ex_cur_inst_addr[9]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_8_ ( .D(n127), .CK(clk), .Q(
        ex_cur_inst_addr[8]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_7_ ( .D(n126), .CK(clk), .Q(
        ex_cur_inst_addr[7]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_6_ ( .D(n125), .CK(clk), .Q(
        ex_cur_inst_addr[6]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_5_ ( .D(n124), .CK(clk), .Q(
        ex_cur_inst_addr[5]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_4_ ( .D(n123), .CK(clk), .Q(
        ex_cur_inst_addr[4]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_3_ ( .D(n122), .CK(clk), .Q(
        ex_cur_inst_addr[3]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_2_ ( .D(n121), .CK(clk), .Q(
        ex_cur_inst_addr[2]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_1_ ( .D(n120), .CK(clk), .Q(
        ex_cur_inst_addr[1]) );
  DQV4_8TH40 ex_cur_inst_addr_reg_0_ ( .D(n119), .CK(clk), .Q(
        ex_cur_inst_addr[0]) );
  DQV4_8TH40 ex_inst_type_reg_7_ ( .D(n118), .CK(clk), .Q(ex_inst_type[7]) );
  DQV4_8TH40 ex_inst_type_reg_6_ ( .D(n117), .CK(clk), .Q(ex_inst_type[6]) );
  DQV4_8TH40 ex_inst_type_reg_5_ ( .D(n116), .CK(clk), .Q(ex_inst_type[5]) );
  DQV4_8TH40 ex_inst_type_reg_4_ ( .D(n115), .CK(clk), .Q(ex_inst_type[4]) );
  DQV4_8TH40 ex_inst_type_reg_3_ ( .D(n114), .CK(clk), .Q(ex_inst_type[3]) );
  DQV4_8TH40 ex_inst_type_reg_2_ ( .D(n113), .CK(clk), .Q(ex_inst_type[2]) );
  DQV4_8TH40 ex_inst_type_reg_1_ ( .D(n112), .CK(clk), .Q(ex_inst_type[1]) );
  DQV4_8TH40 ex_inst_type_reg_0_ ( .D(n111), .CK(clk), .Q(ex_inst_type[0]) );
  DQV4_8TH40 ex_inst_class_reg_2_ ( .D(n110), .CK(clk), .Q(ex_inst_class[2])
         );
  DQV4_8TH40 ex_inst_class_reg_1_ ( .D(n109), .CK(clk), .Q(ex_inst_class[1])
         );
  DQV4_8TH40 ex_inst_class_reg_0_ ( .D(n108), .CK(clk), .Q(ex_inst_class[0])
         );
  DQV4_8TH40 ex_gpr1_data_reg_31_ ( .D(n107), .CK(clk), .Q(ex_gpr1_data[31])
         );
  DQV4_8TH40 ex_gpr1_data_reg_30_ ( .D(n106), .CK(clk), .Q(ex_gpr1_data[30])
         );
  DQV4_8TH40 ex_gpr1_data_reg_29_ ( .D(n105), .CK(clk), .Q(ex_gpr1_data[29])
         );
  DQV4_8TH40 ex_gpr1_data_reg_28_ ( .D(n104), .CK(clk), .Q(ex_gpr1_data[28])
         );
  DQV4_8TH40 ex_gpr1_data_reg_27_ ( .D(n103), .CK(clk), .Q(ex_gpr1_data[27])
         );
  DQV4_8TH40 ex_gpr1_data_reg_26_ ( .D(n102), .CK(clk), .Q(ex_gpr1_data[26])
         );
  DQV4_8TH40 ex_gpr1_data_reg_25_ ( .D(n101), .CK(clk), .Q(ex_gpr1_data[25])
         );
  DQV4_8TH40 ex_gpr1_data_reg_24_ ( .D(n100), .CK(clk), .Q(ex_gpr1_data[24])
         );
  DQV4_8TH40 ex_gpr1_data_reg_23_ ( .D(n99), .CK(clk), .Q(ex_gpr1_data[23]) );
  DQV4_8TH40 ex_gpr1_data_reg_22_ ( .D(n98), .CK(clk), .Q(ex_gpr1_data[22]) );
  DQV4_8TH40 ex_gpr1_data_reg_21_ ( .D(n97), .CK(clk), .Q(ex_gpr1_data[21]) );
  DQV4_8TH40 ex_gpr1_data_reg_20_ ( .D(n96), .CK(clk), .Q(ex_gpr1_data[20]) );
  DQV4_8TH40 ex_gpr1_data_reg_19_ ( .D(n95), .CK(clk), .Q(ex_gpr1_data[19]) );
  DQV4_8TH40 ex_gpr1_data_reg_18_ ( .D(n94), .CK(clk), .Q(ex_gpr1_data[18]) );
  DQV4_8TH40 ex_gpr1_data_reg_17_ ( .D(n93), .CK(clk), .Q(ex_gpr1_data[17]) );
  DQV4_8TH40 ex_gpr1_data_reg_16_ ( .D(n92), .CK(clk), .Q(ex_gpr1_data[16]) );
  DQV4_8TH40 ex_gpr1_data_reg_15_ ( .D(n91), .CK(clk), .Q(ex_gpr1_data[15]) );
  DQV4_8TH40 ex_gpr1_data_reg_14_ ( .D(n90), .CK(clk), .Q(ex_gpr1_data[14]) );
  DQV4_8TH40 ex_gpr1_data_reg_13_ ( .D(n89), .CK(clk), .Q(ex_gpr1_data[13]) );
  DQV4_8TH40 ex_gpr1_data_reg_12_ ( .D(n88), .CK(clk), .Q(ex_gpr1_data[12]) );
  DQV4_8TH40 ex_gpr1_data_reg_11_ ( .D(n87), .CK(clk), .Q(ex_gpr1_data[11]) );
  DQV4_8TH40 ex_gpr1_data_reg_10_ ( .D(n86), .CK(clk), .Q(ex_gpr1_data[10]) );
  DQV4_8TH40 ex_gpr1_data_reg_9_ ( .D(n85), .CK(clk), .Q(ex_gpr1_data[9]) );
  DQV4_8TH40 ex_gpr1_data_reg_8_ ( .D(n84), .CK(clk), .Q(ex_gpr1_data[8]) );
  DQV4_8TH40 ex_gpr1_data_reg_7_ ( .D(n83), .CK(clk), .Q(ex_gpr1_data[7]) );
  DQV4_8TH40 ex_gpr1_data_reg_6_ ( .D(n82), .CK(clk), .Q(ex_gpr1_data[6]) );
  DQV4_8TH40 ex_gpr1_data_reg_5_ ( .D(n81), .CK(clk), .Q(ex_gpr1_data[5]) );
  DQV4_8TH40 ex_gpr1_data_reg_4_ ( .D(n80), .CK(clk), .Q(ex_gpr1_data[4]) );
  DQV4_8TH40 ex_gpr1_data_reg_3_ ( .D(n79), .CK(clk), .Q(ex_gpr1_data[3]) );
  DQV4_8TH40 ex_gpr1_data_reg_2_ ( .D(n78), .CK(clk), .Q(ex_gpr1_data[2]) );
  DQV4_8TH40 ex_gpr1_data_reg_1_ ( .D(n77), .CK(clk), .Q(ex_gpr1_data[1]) );
  DQV4_8TH40 ex_gpr1_data_reg_0_ ( .D(n76), .CK(clk), .Q(ex_gpr1_data[0]) );
  DQV4_8TH40 ex_gpr2_data_reg_31_ ( .D(n75), .CK(clk), .Q(ex_gpr2_data[31]) );
  DQV4_8TH40 ex_gpr2_data_reg_30_ ( .D(n74), .CK(clk), .Q(ex_gpr2_data[30]) );
  DQV4_8TH40 ex_gpr2_data_reg_29_ ( .D(n73), .CK(clk), .Q(ex_gpr2_data[29]) );
  DQV4_8TH40 ex_gpr2_data_reg_28_ ( .D(n72), .CK(clk), .Q(ex_gpr2_data[28]) );
  DQV4_8TH40 ex_gpr2_data_reg_27_ ( .D(n71), .CK(clk), .Q(ex_gpr2_data[27]) );
  DQV4_8TH40 ex_gpr2_data_reg_26_ ( .D(n70), .CK(clk), .Q(ex_gpr2_data[26]) );
  DQV4_8TH40 ex_gpr2_data_reg_25_ ( .D(n69), .CK(clk), .Q(ex_gpr2_data[25]) );
  DQV4_8TH40 ex_gpr2_data_reg_24_ ( .D(n68), .CK(clk), .Q(ex_gpr2_data[24]) );
  DQV4_8TH40 ex_gpr2_data_reg_23_ ( .D(n67), .CK(clk), .Q(ex_gpr2_data[23]) );
  DQV4_8TH40 ex_gpr2_data_reg_22_ ( .D(n66), .CK(clk), .Q(ex_gpr2_data[22]) );
  DQV4_8TH40 ex_gpr2_data_reg_21_ ( .D(n65), .CK(clk), .Q(ex_gpr2_data[21]) );
  DQV4_8TH40 ex_gpr2_data_reg_20_ ( .D(n64), .CK(clk), .Q(ex_gpr2_data[20]) );
  DQV4_8TH40 ex_gpr2_data_reg_19_ ( .D(n63), .CK(clk), .Q(ex_gpr2_data[19]) );
  DQV4_8TH40 ex_gpr2_data_reg_18_ ( .D(n62), .CK(clk), .Q(ex_gpr2_data[18]) );
  DQV4_8TH40 ex_gpr2_data_reg_17_ ( .D(n61), .CK(clk), .Q(ex_gpr2_data[17]) );
  DQV4_8TH40 ex_gpr2_data_reg_16_ ( .D(n60), .CK(clk), .Q(ex_gpr2_data[16]) );
  DQV4_8TH40 ex_gpr2_data_reg_15_ ( .D(n59), .CK(clk), .Q(ex_gpr2_data[15]) );
  DQV4_8TH40 ex_gpr2_data_reg_14_ ( .D(n58), .CK(clk), .Q(ex_gpr2_data[14]) );
  DQV4_8TH40 ex_gpr2_data_reg_13_ ( .D(n57), .CK(clk), .Q(ex_gpr2_data[13]) );
  DQV4_8TH40 ex_gpr2_data_reg_12_ ( .D(n56), .CK(clk), .Q(ex_gpr2_data[12]) );
  DQV4_8TH40 ex_gpr2_data_reg_11_ ( .D(n55), .CK(clk), .Q(ex_gpr2_data[11]) );
  DQV4_8TH40 ex_gpr2_data_reg_10_ ( .D(n54), .CK(clk), .Q(ex_gpr2_data[10]) );
  DQV4_8TH40 ex_gpr2_data_reg_9_ ( .D(n53), .CK(clk), .Q(ex_gpr2_data[9]) );
  DQV4_8TH40 ex_gpr2_data_reg_8_ ( .D(n52), .CK(clk), .Q(ex_gpr2_data[8]) );
  DQV4_8TH40 ex_gpr2_data_reg_7_ ( .D(n51), .CK(clk), .Q(ex_gpr2_data[7]) );
  DQV4_8TH40 ex_gpr2_data_reg_6_ ( .D(n50), .CK(clk), .Q(ex_gpr2_data[6]) );
  DQV4_8TH40 ex_gpr2_data_reg_5_ ( .D(n49), .CK(clk), .Q(ex_gpr2_data[5]) );
  DQV4_8TH40 ex_gpr2_data_reg_4_ ( .D(n48), .CK(clk), .Q(ex_gpr2_data[4]) );
  DQV4_8TH40 ex_gpr2_data_reg_3_ ( .D(n47), .CK(clk), .Q(ex_gpr2_data[3]) );
  DQV4_8TH40 ex_gpr2_data_reg_2_ ( .D(n46), .CK(clk), .Q(ex_gpr2_data[2]) );
  DQV4_8TH40 ex_gpr2_data_reg_1_ ( .D(n45), .CK(clk), .Q(ex_gpr2_data[1]) );
  DQV4_8TH40 ex_gpr2_data_reg_0_ ( .D(n44), .CK(clk), .Q(ex_gpr2_data[0]) );
  DQV4_8TH40 ex_target_gpr_reg_4_ ( .D(n43), .CK(clk), .Q(ex_target_gpr[4]) );
  DQV4_8TH40 ex_target_gpr_reg_3_ ( .D(n42), .CK(clk), .Q(ex_target_gpr[3]) );
  DQV4_8TH40 ex_target_gpr_reg_2_ ( .D(n41), .CK(clk), .Q(ex_target_gpr[2]) );
  DQV4_8TH40 ex_target_gpr_reg_1_ ( .D(n40), .CK(clk), .Q(ex_target_gpr[1]) );
  DQV4_8TH40 ex_target_gpr_reg_0_ ( .D(n39), .CK(clk), .Q(ex_target_gpr[0]) );
  DQV4_8TH40 ex_gpr_we_reg ( .D(n38), .CK(clk), .Q(ex_gpr_we) );
  DQV4_8TH40 ex_link_addr_reg_31_ ( .D(n37), .CK(clk), .Q(ex_link_addr[31]) );
  DQV4_8TH40 ex_link_addr_reg_30_ ( .D(n36), .CK(clk), .Q(ex_link_addr[30]) );
  DQV4_8TH40 ex_link_addr_reg_29_ ( .D(n35), .CK(clk), .Q(ex_link_addr[29]) );
  DQV4_8TH40 ex_link_addr_reg_28_ ( .D(n34), .CK(clk), .Q(ex_link_addr[28]) );
  DQV4_8TH40 ex_link_addr_reg_27_ ( .D(n33), .CK(clk), .Q(ex_link_addr[27]) );
  DQV4_8TH40 ex_link_addr_reg_26_ ( .D(n32), .CK(clk), .Q(ex_link_addr[26]) );
  DQV4_8TH40 ex_link_addr_reg_25_ ( .D(n31), .CK(clk), .Q(ex_link_addr[25]) );
  DQV4_8TH40 ex_link_addr_reg_24_ ( .D(n30), .CK(clk), .Q(ex_link_addr[24]) );
  DQV4_8TH40 ex_link_addr_reg_23_ ( .D(n29), .CK(clk), .Q(ex_link_addr[23]) );
  DQV4_8TH40 ex_link_addr_reg_22_ ( .D(n28), .CK(clk), .Q(ex_link_addr[22]) );
  DQV4_8TH40 ex_link_addr_reg_21_ ( .D(n27), .CK(clk), .Q(ex_link_addr[21]) );
  DQV4_8TH40 ex_link_addr_reg_20_ ( .D(n26), .CK(clk), .Q(ex_link_addr[20]) );
  DQV4_8TH40 ex_link_addr_reg_19_ ( .D(n25), .CK(clk), .Q(ex_link_addr[19]) );
  DQV4_8TH40 ex_link_addr_reg_18_ ( .D(n24), .CK(clk), .Q(ex_link_addr[18]) );
  DQV4_8TH40 ex_link_addr_reg_17_ ( .D(n23), .CK(clk), .Q(ex_link_addr[17]) );
  DQV4_8TH40 ex_link_addr_reg_16_ ( .D(n22), .CK(clk), .Q(ex_link_addr[16]) );
  DQV4_8TH40 ex_link_addr_reg_15_ ( .D(n21), .CK(clk), .Q(ex_link_addr[15]) );
  DQV4_8TH40 ex_link_addr_reg_14_ ( .D(n20), .CK(clk), .Q(ex_link_addr[14]) );
  DQV4_8TH40 ex_link_addr_reg_13_ ( .D(n19), .CK(clk), .Q(ex_link_addr[13]) );
  DQV4_8TH40 ex_link_addr_reg_12_ ( .D(n18), .CK(clk), .Q(ex_link_addr[12]) );
  DQV4_8TH40 ex_link_addr_reg_11_ ( .D(n17), .CK(clk), .Q(ex_link_addr[11]) );
  DQV4_8TH40 ex_link_addr_reg_10_ ( .D(n16), .CK(clk), .Q(ex_link_addr[10]) );
  DQV4_8TH40 ex_link_addr_reg_9_ ( .D(n15), .CK(clk), .Q(ex_link_addr[9]) );
  DQV4_8TH40 ex_link_addr_reg_8_ ( .D(n14), .CK(clk), .Q(ex_link_addr[8]) );
  DQV4_8TH40 ex_link_addr_reg_7_ ( .D(n13), .CK(clk), .Q(ex_link_addr[7]) );
  DQV4_8TH40 ex_link_addr_reg_6_ ( .D(n12), .CK(clk), .Q(ex_link_addr[6]) );
  DQV4_8TH40 ex_link_addr_reg_5_ ( .D(n11), .CK(clk), .Q(ex_link_addr[5]) );
  DQV4_8TH40 ex_link_addr_reg_4_ ( .D(n10), .CK(clk), .Q(ex_link_addr[4]) );
  DQV4_8TH40 ex_link_addr_reg_3_ ( .D(n9), .CK(clk), .Q(ex_link_addr[3]) );
  DQV4_8TH40 ex_link_addr_reg_2_ ( .D(n8), .CK(clk), .Q(ex_link_addr[2]) );
  DQV4_8TH40 ex_link_addr_reg_1_ ( .D(n7), .CK(clk), .Q(ex_link_addr[1]) );
  DQV4_8TH40 ex_link_addr_reg_0_ ( .D(n6), .CK(clk), .Q(ex_link_addr[0]) );
  DQV4_8TH40 ex_inst_delayslot_reg ( .D(n5), .CK(clk), .Q(ex_inst_delayslot)
         );
  DQV4_8TH40 nxt_inst_delayslot_reg ( .D(n4), .CK(clk), .Q(nxt_inst_delayslot)
         );
  CLKBUFV2_8TH40 U2 ( .I(n175), .Z(n169) );
  CLKBUFV2_8TH40 U3 ( .I(n161), .Z(n154) );
  AO22V4_8TH40 U4 ( .A1(ex_inst_type[1]), .A2(n151), .B1(id_inst_type[1]), 
        .B2(n162), .Z(n112) );
  AO22V4_8TH40 U5 ( .A1(ex_link_addr[5]), .A2(n152), .B1(id_link_addr[5]), 
        .B2(n164), .Z(n11) );
  AO22V4_8TH40 U6 ( .A1(ex_link_addr[6]), .A2(n2), .B1(id_link_addr[6]), .B2(
        n162), .Z(n12) );
  AO22V4_8TH40 U7 ( .A1(ex_link_addr[7]), .A2(n177), .B1(id_link_addr[7]), 
        .B2(n178), .Z(n13) );
  AO22V4_8TH40 U8 ( .A1(ex_link_addr[8]), .A2(n152), .B1(id_link_addr[8]), 
        .B2(n178), .Z(n14) );
  AO22V4_8TH40 U9 ( .A1(ex_link_addr[9]), .A2(n177), .B1(id_link_addr[9]), 
        .B2(n164), .Z(n15) );
  AO22V4_8TH40 U10 ( .A1(ex_link_addr[10]), .A2(n153), .B1(id_link_addr[10]), 
        .B2(n164), .Z(n16) );
  AO22V4_8TH40 U11 ( .A1(ex_link_addr[11]), .A2(n151), .B1(id_link_addr[11]), 
        .B2(n165), .Z(n17) );
  AO22V4_8TH40 U12 ( .A1(ex_link_addr[12]), .A2(n3), .B1(id_link_addr[12]), 
        .B2(n165), .Z(n18) );
  AO22V4_8TH40 U13 ( .A1(ex_link_addr[13]), .A2(n177), .B1(id_link_addr[13]), 
        .B2(n165), .Z(n19) );
  AO22V4_8TH40 U14 ( .A1(ex_link_addr[14]), .A2(n151), .B1(id_link_addr[14]), 
        .B2(n166), .Z(n20) );
  AO22V4_8TH40 U15 ( .A1(ex_link_addr[15]), .A2(n151), .B1(id_link_addr[15]), 
        .B2(n166), .Z(n21) );
  AO22V4_8TH40 U16 ( .A1(ex_link_addr[16]), .A2(n151), .B1(id_link_addr[16]), 
        .B2(n166), .Z(n22) );
  AO22V4_8TH40 U17 ( .A1(ex_link_addr[17]), .A2(n151), .B1(id_link_addr[17]), 
        .B2(n166), .Z(n23) );
  AO22V4_8TH40 U18 ( .A1(ex_link_addr[18]), .A2(n151), .B1(id_link_addr[18]), 
        .B2(n164), .Z(n24) );
  AO22V4_8TH40 U19 ( .A1(ex_link_addr[19]), .A2(n151), .B1(id_link_addr[19]), 
        .B2(n165), .Z(n25) );
  AO22V4_8TH40 U20 ( .A1(ex_link_addr[20]), .A2(n151), .B1(id_link_addr[20]), 
        .B2(n166), .Z(n26) );
  AO22V4_8TH40 U21 ( .A1(ex_link_addr[21]), .A2(n151), .B1(id_link_addr[21]), 
        .B2(n168), .Z(n27) );
  AO22V4_8TH40 U22 ( .A1(ex_link_addr[22]), .A2(n151), .B1(id_link_addr[22]), 
        .B2(n176), .Z(n28) );
  AO22V4_8TH40 U23 ( .A1(ex_link_addr[23]), .A2(n152), .B1(id_link_addr[23]), 
        .B2(n167), .Z(n29) );
  AO22V4_8TH40 U24 ( .A1(ex_link_addr[24]), .A2(n3), .B1(id_link_addr[24]), 
        .B2(n162), .Z(n30) );
  AO22V4_8TH40 U25 ( .A1(ex_link_addr[25]), .A2(n177), .B1(id_link_addr[25]), 
        .B2(n178), .Z(n31) );
  AO22V4_8TH40 U26 ( .A1(ex_link_addr[26]), .A2(n153), .B1(id_link_addr[26]), 
        .B2(n164), .Z(n32) );
  AO22V4_8TH40 U27 ( .A1(ex_link_addr[27]), .A2(n2), .B1(id_link_addr[27]), 
        .B2(n165), .Z(n33) );
  AO22V4_8TH40 U28 ( .A1(ex_link_addr[28]), .A2(n1), .B1(id_link_addr[28]), 
        .B2(n166), .Z(n34) );
  AO22V4_8TH40 U29 ( .A1(ex_link_addr[29]), .A2(n151), .B1(id_link_addr[29]), 
        .B2(n168), .Z(n35) );
  AO22V4_8TH40 U30 ( .A1(ex_link_addr[30]), .A2(n152), .B1(id_link_addr[30]), 
        .B2(n167), .Z(n36) );
  AO22V4_8TH40 U31 ( .A1(ex_gpr_we), .A2(n3), .B1(id_gpr_we), .B2(n167), .Z(
        n38) );
  AO22V4_8TH40 U32 ( .A1(ex_inst_type[4]), .A2(n1), .B1(id_inst_type[4]), .B2(
        n162), .Z(n115) );
  AO22V4_8TH40 U33 ( .A1(ex_inst_type[0]), .A2(n1), .B1(id_inst_type[0]), .B2(
        n162), .Z(n111) );
  AO22V4_8TH40 U34 ( .A1(ex_inst_type[2]), .A2(n177), .B1(id_inst_type[2]), 
        .B2(n162), .Z(n113) );
  AO22V4_8TH40 U35 ( .A1(ex_inst_type[3]), .A2(n153), .B1(id_inst_type[3]), 
        .B2(n162), .Z(n114) );
  AO22V4_8TH40 U36 ( .A1(ex_inst_type[5]), .A2(n177), .B1(id_inst_type[5]), 
        .B2(n162), .Z(n116) );
  AO22V4_8TH40 U37 ( .A1(ex_except_type[9]), .A2(n152), .B1(id_except_type[9]), 
        .B2(n164), .Z(n160) );
  AO22V4_8TH40 U38 ( .A1(ex_link_addr[0]), .A2(n177), .B1(id_link_addr[0]), 
        .B2(n168), .Z(n6) );
  AO22V4_8TH40 U39 ( .A1(ex_link_addr[1]), .A2(n2), .B1(id_link_addr[1]), .B2(
        n167), .Z(n7) );
  AO22V4_8TH40 U40 ( .A1(ex_link_addr[2]), .A2(n1), .B1(id_link_addr[2]), .B2(
        n168), .Z(n8) );
  AO22V4_8TH40 U41 ( .A1(ex_target_gpr[0]), .A2(n177), .B1(id_target_gpr[0]), 
        .B2(n167), .Z(n39) );
  AO22V4_8TH40 U42 ( .A1(ex_target_gpr[1]), .A2(n3), .B1(id_target_gpr[1]), 
        .B2(n167), .Z(n40) );
  AO22V4_8TH40 U43 ( .A1(ex_target_gpr[2]), .A2(n3), .B1(id_target_gpr[2]), 
        .B2(n167), .Z(n41) );
  AO22V4_8TH40 U44 ( .A1(ex_target_gpr[3]), .A2(n3), .B1(id_target_gpr[3]), 
        .B2(n167), .Z(n42) );
  AO22V4_8TH40 U45 ( .A1(ex_target_gpr[4]), .A2(n3), .B1(id_target_gpr[4]), 
        .B2(n167), .Z(n43) );
  AO22V4_8TH40 U46 ( .A1(ex_inst_class[1]), .A2(n3), .B1(id_inst_class[1]), 
        .B2(n165), .Z(n109) );
  AO22V4_8TH40 U47 ( .A1(ex_inst_class[2]), .A2(n151), .B1(id_inst_class[2]), 
        .B2(n162), .Z(n110) );
  AO22V4_8TH40 U48 ( .A1(ex_inst_type[6]), .A2(n152), .B1(id_inst_type[6]), 
        .B2(n162), .Z(n117) );
  AO22V4_8TH40 U49 ( .A1(ex_except_type[12]), .A2(n2), .B1(id_except_type[12]), 
        .B2(n165), .Z(n163) );
  AO22V4_8TH40 U50 ( .A1(ex_link_addr[4]), .A2(n153), .B1(id_link_addr[4]), 
        .B2(n166), .Z(n10) );
  AO22V4_8TH40 U51 ( .A1(ex_inst_class[0]), .A2(n153), .B1(id_inst_class[0]), 
        .B2(n176), .Z(n108) );
  AO22V4_8TH40 U52 ( .A1(ex_link_addr[3]), .A2(n153), .B1(id_link_addr[3]), 
        .B2(n168), .Z(n9) );
  AO22V4_8TH40 U53 ( .A1(ex_inst_delayslot), .A2(n3), .B1(id_inst_delayslot), 
        .B2(n176), .Z(n5) );
  AO22V4_8TH40 U54 ( .A1(ex_link_addr[31]), .A2(n153), .B1(id_link_addr[31]), 
        .B2(n167), .Z(n37) );
  AO22V4_8TH40 U55 ( .A1(ex_except_type[8]), .A2(n1), .B1(id_except_type[8]), 
        .B2(n164), .Z(n159) );
  AND4V2_8TH40 U56 ( .A1(n180), .A2(flush_BAR), .A3(stall_ctrl[2]), .A4(n179), 
        .Z(n177) );
  INV2_8TH40 U57 ( .I(n170), .ZN(n167) );
  INV2_8TH40 U58 ( .I(n171), .ZN(n166) );
  CLKBUFV2_8TH40 U59 ( .I(n175), .Z(n170) );
  CLKBUFV2_8TH40 U60 ( .I(n173), .Z(n171) );
  INV2_8TH40 U61 ( .I(n157), .ZN(n3) );
  INV2_8TH40 U62 ( .I(n158), .ZN(n2) );
  INV2_8TH40 U63 ( .I(n158), .ZN(n1) );
  INV2_8TH40 U64 ( .I(n155), .ZN(n152) );
  INV2_8TH40 U65 ( .I(n156), .ZN(n151) );
  INV2_8TH40 U66 ( .I(n169), .ZN(n168) );
  INV2_8TH40 U67 ( .I(n173), .ZN(n162) );
  INV2_8TH40 U68 ( .I(n172), .ZN(n164) );
  INV2_8TH40 U69 ( .I(n172), .ZN(n165) );
  CLKBUFV2_8TH40 U70 ( .I(n155), .Z(n157) );
  CLKBUFV2_8TH40 U71 ( .I(n156), .Z(n158) );
  CLKBUFV2_8TH40 U72 ( .I(n161), .Z(n155) );
  CLKBUFV2_8TH40 U73 ( .I(n161), .Z(n156) );
  CLKBUFV2_8TH40 U74 ( .I(n174), .Z(n173) );
  CLKBUFV2_8TH40 U75 ( .I(n174), .Z(n172) );
  INV2_8TH40 U76 ( .I(n176), .ZN(n175) );
  INV2_8TH40 U77 ( .I(n154), .ZN(n153) );
  CLKBUFV2_8TH40 U78 ( .I(n178), .Z(n176) );
  INV2_8TH40 U79 ( .I(n177), .ZN(n161) );
  INV2_8TH40 U80 ( .I(n178), .ZN(n174) );
  AO22V0_8TH40 U81 ( .A1(ex_gpr1_data[23]), .A2(n2), .B1(id_gpr1_data[23]), 
        .B2(n176), .Z(n99) );
  AO22V0_8TH40 U82 ( .A1(ex_gpr1_data[22]), .A2(n153), .B1(id_gpr1_data[22]), 
        .B2(n176), .Z(n98) );
  AO22V0_8TH40 U83 ( .A1(ex_gpr1_data[21]), .A2(n177), .B1(id_gpr1_data[21]), 
        .B2(n178), .Z(n97) );
  AO22V0_8TH40 U84 ( .A1(ex_gpr1_data[20]), .A2(n3), .B1(id_gpr1_data[20]), 
        .B2(n176), .Z(n96) );
  AO22V0_8TH40 U85 ( .A1(ex_gpr1_data[19]), .A2(n152), .B1(id_gpr1_data[19]), 
        .B2(n178), .Z(n95) );
  AO22V0_8TH40 U86 ( .A1(ex_gpr1_data[18]), .A2(n151), .B1(id_gpr1_data[18]), 
        .B2(n176), .Z(n94) );
  AO22V0_8TH40 U87 ( .A1(ex_gpr1_data[17]), .A2(n1), .B1(id_gpr1_data[17]), 
        .B2(n178), .Z(n93) );
  AO22V0_8TH40 U88 ( .A1(ex_gpr1_data[16]), .A2(n1), .B1(id_gpr1_data[16]), 
        .B2(n176), .Z(n92) );
  AO22V0_8TH40 U89 ( .A1(ex_gpr1_data[15]), .A2(n2), .B1(id_gpr1_data[15]), 
        .B2(n178), .Z(n91) );
  AO22V0_8TH40 U90 ( .A1(ex_gpr1_data[14]), .A2(n153), .B1(id_gpr1_data[14]), 
        .B2(n176), .Z(n90) );
  AO22V0_8TH40 U91 ( .A1(ex_gpr1_data[13]), .A2(n177), .B1(id_gpr1_data[13]), 
        .B2(n168), .Z(n89) );
  AO22V0_8TH40 U92 ( .A1(ex_gpr1_data[12]), .A2(n3), .B1(id_gpr1_data[12]), 
        .B2(n168), .Z(n88) );
  AO22V0_8TH40 U93 ( .A1(ex_gpr1_data[11]), .A2(n1), .B1(id_gpr1_data[11]), 
        .B2(n168), .Z(n87) );
  AO22V0_8TH40 U94 ( .A1(ex_gpr1_data[10]), .A2(n1), .B1(id_gpr1_data[10]), 
        .B2(n168), .Z(n86) );
  AO22V0_8TH40 U95 ( .A1(ex_gpr1_data[9]), .A2(n1), .B1(id_gpr1_data[9]), .B2(
        n168), .Z(n85) );
  AO22V0_8TH40 U96 ( .A1(ex_gpr1_data[8]), .A2(n1), .B1(id_gpr1_data[8]), .B2(
        n168), .Z(n84) );
  AO22V0_8TH40 U97 ( .A1(ex_gpr1_data[7]), .A2(n1), .B1(id_gpr1_data[7]), .B2(
        n168), .Z(n83) );
  AO22V0_8TH40 U98 ( .A1(ex_gpr1_data[6]), .A2(n1), .B1(id_gpr1_data[6]), .B2(
        n168), .Z(n82) );
  AO22V0_8TH40 U99 ( .A1(ex_gpr1_data[5]), .A2(n1), .B1(id_gpr1_data[5]), .B2(
        n168), .Z(n81) );
  AO22V0_8TH40 U100 ( .A1(ex_gpr1_data[4]), .A2(n1), .B1(id_gpr1_data[4]), 
        .B2(n168), .Z(n80) );
  AO22V0_8TH40 U101 ( .A1(ex_gpr1_data[3]), .A2(n1), .B1(id_gpr1_data[3]), 
        .B2(n167), .Z(n79) );
  AO22V0_8TH40 U102 ( .A1(ex_gpr1_data[2]), .A2(n1), .B1(id_gpr1_data[2]), 
        .B2(n166), .Z(n78) );
  AO22V0_8TH40 U103 ( .A1(ex_gpr1_data[1]), .A2(n1), .B1(id_gpr1_data[1]), 
        .B2(n168), .Z(n77) );
  AO22V0_8TH40 U104 ( .A1(ex_gpr1_data[0]), .A2(n1), .B1(id_gpr1_data[0]), 
        .B2(n164), .Z(n76) );
  AO22V0_8TH40 U105 ( .A1(ex_gpr2_data[31]), .A2(n2), .B1(id_gpr2_data[31]), 
        .B2(n165), .Z(n75) );
  AO22V0_8TH40 U106 ( .A1(ex_gpr2_data[30]), .A2(n2), .B1(id_gpr2_data[30]), 
        .B2(n176), .Z(n74) );
  AO22V0_8TH40 U107 ( .A1(ex_gpr2_data[29]), .A2(n2), .B1(id_gpr2_data[29]), 
        .B2(n168), .Z(n73) );
  AO22V0_8TH40 U108 ( .A1(ex_gpr2_data[28]), .A2(n2), .B1(id_gpr2_data[28]), 
        .B2(n162), .Z(n72) );
  AO22V0_8TH40 U109 ( .A1(ex_gpr2_data[27]), .A2(n2), .B1(id_gpr2_data[27]), 
        .B2(n167), .Z(n71) );
  AO22V0_8TH40 U110 ( .A1(ex_gpr2_data[26]), .A2(n2), .B1(id_gpr2_data[26]), 
        .B2(n178), .Z(n70) );
  AO22V0_8TH40 U111 ( .A1(ex_gpr2_data[25]), .A2(n2), .B1(id_gpr2_data[25]), 
        .B2(n162), .Z(n69) );
  AO22V0_8TH40 U112 ( .A1(ex_gpr2_data[24]), .A2(n2), .B1(id_gpr2_data[24]), 
        .B2(n162), .Z(n68) );
  AO22V0_8TH40 U113 ( .A1(ex_gpr2_data[23]), .A2(n2), .B1(id_gpr2_data[23]), 
        .B2(n176), .Z(n67) );
  AO22V0_8TH40 U114 ( .A1(ex_gpr2_data[22]), .A2(n2), .B1(id_gpr2_data[22]), 
        .B2(n168), .Z(n66) );
  AO22V0_8TH40 U115 ( .A1(ex_gpr2_data[21]), .A2(n2), .B1(id_gpr2_data[21]), 
        .B2(n178), .Z(n65) );
  AO22V0_8TH40 U116 ( .A1(ex_gpr2_data[20]), .A2(n2), .B1(id_gpr2_data[20]), 
        .B2(n167), .Z(n64) );
  AO22V0_8TH40 U117 ( .A1(ex_gpr2_data[19]), .A2(n153), .B1(id_gpr2_data[19]), 
        .B2(n178), .Z(n63) );
  AO22V0_8TH40 U118 ( .A1(ex_gpr2_data[18]), .A2(n152), .B1(id_gpr2_data[18]), 
        .B2(n166), .Z(n62) );
  AO22V0_8TH40 U119 ( .A1(ex_gpr2_data[17]), .A2(n1), .B1(id_gpr2_data[17]), 
        .B2(n176), .Z(n61) );
  AO22V0_8TH40 U120 ( .A1(ex_gpr2_data[16]), .A2(n2), .B1(id_gpr2_data[16]), 
        .B2(n164), .Z(n60) );
  AO22V0_8TH40 U121 ( .A1(ex_gpr2_data[15]), .A2(n152), .B1(id_gpr2_data[15]), 
        .B2(n165), .Z(n59) );
  AO22V0_8TH40 U122 ( .A1(ex_gpr2_data[14]), .A2(n177), .B1(id_gpr2_data[14]), 
        .B2(n176), .Z(n58) );
  AO22V0_8TH40 U123 ( .A1(ex_gpr2_data[13]), .A2(n152), .B1(id_gpr2_data[13]), 
        .B2(n165), .Z(n57) );
  AO22V0_8TH40 U124 ( .A1(ex_gpr2_data[12]), .A2(n153), .B1(id_gpr2_data[12]), 
        .B2(n176), .Z(n56) );
  AO22V0_8TH40 U125 ( .A1(ex_gpr2_data[11]), .A2(n152), .B1(id_gpr2_data[11]), 
        .B2(n167), .Z(n55) );
  AO22V0_8TH40 U126 ( .A1(ex_gpr2_data[10]), .A2(n1), .B1(id_gpr2_data[10]), 
        .B2(n168), .Z(n54) );
  AO22V0_8TH40 U127 ( .A1(ex_gpr2_data[9]), .A2(n2), .B1(id_gpr2_data[9]), 
        .B2(n162), .Z(n53) );
  AO22V0_8TH40 U128 ( .A1(ex_gpr2_data[8]), .A2(n151), .B1(id_gpr2_data[8]), 
        .B2(n178), .Z(n52) );
  AO22V0_8TH40 U129 ( .A1(ex_gpr2_data[7]), .A2(n3), .B1(id_gpr2_data[7]), 
        .B2(n178), .Z(n51) );
  AO22V0_8TH40 U130 ( .A1(ex_gpr2_data[6]), .A2(n3), .B1(id_gpr2_data[6]), 
        .B2(n166), .Z(n50) );
  AO22V0_8TH40 U131 ( .A1(ex_gpr2_data[5]), .A2(n3), .B1(id_gpr2_data[5]), 
        .B2(n162), .Z(n49) );
  AO22V0_8TH40 U132 ( .A1(ex_gpr2_data[4]), .A2(n3), .B1(id_gpr2_data[4]), 
        .B2(n164), .Z(n48) );
  AO22V0_8TH40 U133 ( .A1(ex_gpr2_data[3]), .A2(n3), .B1(id_gpr2_data[3]), 
        .B2(n165), .Z(n47) );
  AO22V0_8TH40 U134 ( .A1(ex_gpr2_data[2]), .A2(n3), .B1(id_gpr2_data[2]), 
        .B2(n167), .Z(n46) );
  AO22V0_8TH40 U135 ( .A1(ex_gpr2_data[1]), .A2(n3), .B1(id_gpr2_data[1]), 
        .B2(n167), .Z(n45) );
  AO22V0_8TH40 U136 ( .A1(ex_gpr2_data[0]), .A2(n3), .B1(id_gpr2_data[0]), 
        .B2(n167), .Z(n44) );
  AO22V0_8TH40 U137 ( .A1(nxt_inst_delayslot), .A2(n2), .B1(
        nxtid_inst_delayslot), .B2(n167), .Z(n4) );
  AO22V0_8TH40 U138 ( .A1(ex_inst[15]), .A2(n151), .B1(id_inst[15]), .B2(n166), 
        .Z(n198) );
  AO22V0_8TH40 U139 ( .A1(ex_inst[14]), .A2(n151), .B1(id_inst[14]), .B2(n166), 
        .Z(n197) );
  AO22V0_8TH40 U140 ( .A1(ex_inst[13]), .A2(n151), .B1(id_inst[13]), .B2(n166), 
        .Z(n196) );
  AO22V0_8TH40 U141 ( .A1(ex_inst[12]), .A2(n151), .B1(id_inst[12]), .B2(n166), 
        .Z(n195) );
  AO22V0_8TH40 U142 ( .A1(ex_inst[11]), .A2(n151), .B1(id_inst[11]), .B2(n166), 
        .Z(n194) );
  AO22V0_8TH40 U143 ( .A1(ex_inst[10]), .A2(n3), .B1(id_inst[10]), .B2(n166), 
        .Z(n193) );
  AO22V0_8TH40 U144 ( .A1(ex_inst[9]), .A2(n2), .B1(id_inst[9]), .B2(n166), 
        .Z(n192) );
  AO22V0_8TH40 U145 ( .A1(ex_inst[8]), .A2(n1), .B1(id_inst[8]), .B2(n166), 
        .Z(n191) );
  AO22V0_8TH40 U146 ( .A1(ex_inst[7]), .A2(n2), .B1(id_inst[7]), .B2(n165), 
        .Z(n190) );
  AO22V0_8TH40 U147 ( .A1(ex_inst[6]), .A2(n152), .B1(id_inst[6]), .B2(n165), 
        .Z(n189) );
  AO22V0_8TH40 U148 ( .A1(ex_inst[5]), .A2(n151), .B1(id_inst[5]), .B2(n165), 
        .Z(n188) );
  AO22V0_8TH40 U149 ( .A1(ex_inst[4]), .A2(n153), .B1(id_inst[4]), .B2(n165), 
        .Z(n187) );
  AO22V0_8TH40 U150 ( .A1(ex_inst[3]), .A2(n3), .B1(id_inst[3]), .B2(n165), 
        .Z(n186) );
  AO22V0_8TH40 U151 ( .A1(ex_inst[2]), .A2(n1), .B1(id_inst[2]), .B2(n165), 
        .Z(n185) );
  AO22V0_8TH40 U152 ( .A1(ex_inst[1]), .A2(n1), .B1(id_inst[1]), .B2(n165), 
        .Z(n184) );
  AO22V0_8TH40 U153 ( .A1(ex_inst[0]), .A2(n2), .B1(id_inst[0]), .B2(n165), 
        .Z(n183) );
  AO22V0_8TH40 U154 ( .A1(ex_cur_inst_addr[31]), .A2(n3), .B1(
        id_cur_inst_addr[31]), .B2(n164), .Z(n150) );
  AO22V0_8TH40 U155 ( .A1(ex_cur_inst_addr[30]), .A2(n2), .B1(
        id_cur_inst_addr[30]), .B2(n164), .Z(n149) );
  AO22V0_8TH40 U156 ( .A1(ex_cur_inst_addr[29]), .A2(n153), .B1(
        id_cur_inst_addr[29]), .B2(n164), .Z(n148) );
  AO22V0_8TH40 U157 ( .A1(ex_cur_inst_addr[28]), .A2(n177), .B1(
        id_cur_inst_addr[28]), .B2(n164), .Z(n147) );
  AO22V0_8TH40 U158 ( .A1(ex_cur_inst_addr[27]), .A2(n152), .B1(
        id_cur_inst_addr[27]), .B2(n164), .Z(n146) );
  AO22V0_8TH40 U159 ( .A1(ex_cur_inst_addr[26]), .A2(n2), .B1(
        id_cur_inst_addr[26]), .B2(n164), .Z(n145) );
  AO22V0_8TH40 U160 ( .A1(ex_cur_inst_addr[25]), .A2(n3), .B1(
        id_cur_inst_addr[25]), .B2(n164), .Z(n144) );
  AO22V0_8TH40 U161 ( .A1(ex_cur_inst_addr[24]), .A2(n152), .B1(
        id_cur_inst_addr[24]), .B2(n164), .Z(n143) );
  AO22V0_8TH40 U162 ( .A1(ex_cur_inst_addr[23]), .A2(n152), .B1(
        id_cur_inst_addr[23]), .B2(n166), .Z(n142) );
  AO22V0_8TH40 U163 ( .A1(ex_cur_inst_addr[22]), .A2(n152), .B1(
        id_cur_inst_addr[22]), .B2(n168), .Z(n141) );
  AO22V0_8TH40 U164 ( .A1(ex_cur_inst_addr[21]), .A2(n152), .B1(
        id_cur_inst_addr[21]), .B2(n166), .Z(n140) );
  AO22V0_8TH40 U165 ( .A1(ex_cur_inst_addr[20]), .A2(n152), .B1(
        id_cur_inst_addr[20]), .B2(n178), .Z(n139) );
  AO22V0_8TH40 U166 ( .A1(ex_cur_inst_addr[19]), .A2(n152), .B1(
        id_cur_inst_addr[19]), .B2(n164), .Z(n138) );
  AO22V0_8TH40 U167 ( .A1(ex_cur_inst_addr[18]), .A2(n152), .B1(
        id_cur_inst_addr[18]), .B2(n165), .Z(n137) );
  AO22V0_8TH40 U168 ( .A1(ex_cur_inst_addr[17]), .A2(n152), .B1(
        id_cur_inst_addr[17]), .B2(n176), .Z(n136) );
  AO22V0_8TH40 U169 ( .A1(ex_cur_inst_addr[16]), .A2(n152), .B1(
        id_cur_inst_addr[16]), .B2(n167), .Z(n135) );
  AO22V0_8TH40 U170 ( .A1(ex_cur_inst_addr[15]), .A2(n152), .B1(
        id_cur_inst_addr[15]), .B2(n168), .Z(n134) );
  AO22V0_8TH40 U171 ( .A1(ex_cur_inst_addr[14]), .A2(n152), .B1(
        id_cur_inst_addr[14]), .B2(n162), .Z(n133) );
  AO22V0_8TH40 U172 ( .A1(ex_cur_inst_addr[13]), .A2(n152), .B1(
        id_cur_inst_addr[13]), .B2(n178), .Z(n132) );
  AO22V0_8TH40 U173 ( .A1(ex_cur_inst_addr[12]), .A2(n153), .B1(
        id_cur_inst_addr[12]), .B2(n176), .Z(n131) );
  AO22V0_8TH40 U174 ( .A1(ex_cur_inst_addr[11]), .A2(n177), .B1(
        id_cur_inst_addr[11]), .B2(n178), .Z(n130) );
  AO22V0_8TH40 U175 ( .A1(ex_cur_inst_addr[10]), .A2(n153), .B1(
        id_cur_inst_addr[10]), .B2(n176), .Z(n129) );
  AO22V0_8TH40 U176 ( .A1(ex_cur_inst_addr[9]), .A2(n177), .B1(
        id_cur_inst_addr[9]), .B2(n178), .Z(n128) );
  AO22V0_8TH40 U177 ( .A1(ex_cur_inst_addr[8]), .A2(n177), .B1(
        id_cur_inst_addr[8]), .B2(n176), .Z(n127) );
  AO22V0_8TH40 U178 ( .A1(ex_cur_inst_addr[7]), .A2(n177), .B1(
        id_cur_inst_addr[7]), .B2(n178), .Z(n126) );
  AO22V0_8TH40 U179 ( .A1(ex_cur_inst_addr[6]), .A2(n177), .B1(
        id_cur_inst_addr[6]), .B2(n176), .Z(n125) );
  AO22V0_8TH40 U180 ( .A1(ex_cur_inst_addr[5]), .A2(n177), .B1(
        id_cur_inst_addr[5]), .B2(n178), .Z(n124) );
  AO22V0_8TH40 U181 ( .A1(ex_cur_inst_addr[4]), .A2(n177), .B1(
        id_cur_inst_addr[4]), .B2(n176), .Z(n123) );
  AO22V0_8TH40 U182 ( .A1(ex_cur_inst_addr[3]), .A2(n177), .B1(
        id_cur_inst_addr[3]), .B2(n178), .Z(n122) );
  AO22V0_8TH40 U183 ( .A1(ex_cur_inst_addr[2]), .A2(n177), .B1(
        id_cur_inst_addr[2]), .B2(n164), .Z(n121) );
  AO22V0_8TH40 U184 ( .A1(ex_cur_inst_addr[1]), .A2(n177), .B1(
        id_cur_inst_addr[1]), .B2(n162), .Z(n120) );
  AO22V0_8TH40 U185 ( .A1(ex_cur_inst_addr[0]), .A2(n151), .B1(
        id_cur_inst_addr[0]), .B2(n162), .Z(n119) );
  AO22V0_8TH40 U186 ( .A1(ex_inst_type[7]), .A2(n1), .B1(id_inst_type[7]), 
        .B2(n162), .Z(n118) );
  AO22V0_8TH40 U187 ( .A1(ex_gpr1_data[31]), .A2(n153), .B1(id_gpr1_data[31]), 
        .B2(n164), .Z(n107) );
  AO22V0_8TH40 U188 ( .A1(ex_gpr1_data[30]), .A2(n153), .B1(id_gpr1_data[30]), 
        .B2(n165), .Z(n106) );
  AO22V0_8TH40 U189 ( .A1(ex_gpr1_data[29]), .A2(n153), .B1(id_gpr1_data[29]), 
        .B2(n166), .Z(n105) );
  AO22V0_8TH40 U190 ( .A1(ex_gpr1_data[28]), .A2(n153), .B1(id_gpr1_data[28]), 
        .B2(n168), .Z(n104) );
  AO22V0_8TH40 U191 ( .A1(ex_gpr1_data[27]), .A2(n153), .B1(id_gpr1_data[27]), 
        .B2(n176), .Z(n103) );
  AO22V0_8TH40 U192 ( .A1(ex_gpr1_data[26]), .A2(n153), .B1(id_gpr1_data[26]), 
        .B2(n167), .Z(n102) );
  AO22V0_8TH40 U193 ( .A1(ex_gpr1_data[25]), .A2(n153), .B1(id_gpr1_data[25]), 
        .B2(n162), .Z(n101) );
  AO22V0_8TH40 U194 ( .A1(ex_gpr1_data[24]), .A2(n153), .B1(id_gpr1_data[24]), 
        .B2(n178), .Z(n100) );
  I2NOR4V0_8TH40 U195 ( .A1(flush_BAR), .A2(n179), .B1(n153), .B2(rst), .ZN(
        n178) );
  INAND2V0_8TH40 U196 ( .A1(stall_ctrl[3]), .B1(stall_ctrl[2]), .ZN(n179) );
  CLKNV1_8TH40 U197 ( .I(rst), .ZN(n180) );
endmodule


module inst_execute_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_2__1_,
         ML_int_2__0_, ML_int_3__31_, ML_int_3__30_, ML_int_3__29_,
         ML_int_3__28_, ML_int_3__27_, ML_int_3__26_, ML_int_3__25_,
         ML_int_3__24_, ML_int_3__23_, ML_int_3__22_, ML_int_3__21_,
         ML_int_3__20_, ML_int_3__19_, ML_int_3__18_, ML_int_3__17_,
         ML_int_3__16_, ML_int_3__15_, ML_int_3__14_, ML_int_3__13_,
         ML_int_3__12_, ML_int_3__11_, ML_int_3__10_, ML_int_3__9_,
         ML_int_3__8_, ML_int_3__7_, ML_int_3__6_, ML_int_3__5_, ML_int_3__4_,
         ML_int_3__3_, ML_int_3__2_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__15_,
         ML_int_4__14_, ML_int_4__13_, ML_int_4__12_, ML_int_4__11_,
         ML_int_4__10_, ML_int_4__9_, ML_int_4__8_, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  CKMUX2V4_8TH40 M1_4_30 ( .I0(ML_int_4__30_), .I1(ML_int_4__14_), .S(SH[4]), 
        .Z(B[30]) );
  CKMUX2V4_8TH40 M1_4_28 ( .I0(ML_int_4__28_), .I1(ML_int_4__12_), .S(SH[4]), 
        .Z(B[28]) );
  CKMUX2V4_8TH40 M1_3_31 ( .I0(ML_int_3__31_), .I1(ML_int_3__23_), .S(SH[3]), 
        .Z(ML_int_4__31_) );
  CKMUX2V4_8TH40 M1_3_29 ( .I0(ML_int_3__29_), .I1(ML_int_3__21_), .S(SH[3]), 
        .Z(ML_int_4__29_) );
  CKMUX2V4_8TH40 M1_2_30 ( .I0(ML_int_2__30_), .I1(ML_int_2__26_), .S(SH[2]), 
        .Z(ML_int_3__30_) );
  CKMUX2V2_8TH40 M1_0_31 ( .I0(A[31]), .I1(A[30]), .S(SH[0]), .Z(ML_int_1__31_) );
  CKMUX2V2_8TH40 M1_0_30 ( .I0(A[30]), .I1(A[29]), .S(SH[0]), .Z(ML_int_1__30_) );
  CKMUX2V2_8TH40 M1_1_28 ( .I0(ML_int_1__28_), .I1(ML_int_1__26_), .S(SH[1]), 
        .Z(ML_int_2__28_) );
  CKMUX2V2_8TH40 M1_1_29 ( .I0(ML_int_1__29_), .I1(ML_int_1__27_), .S(SH[1]), 
        .Z(ML_int_2__29_) );
  CKMUX2V2_8TH40 M1_3_15 ( .I0(ML_int_3__15_), .I1(ML_int_3__7_), .S(SH[3]), 
        .Z(ML_int_4__15_) );
  CKMUX2V2_8TH40 M1_3_13 ( .I0(ML_int_3__13_), .I1(ML_int_3__5_), .S(SH[3]), 
        .Z(ML_int_4__13_) );
  CKMUX2V2_8TH40 M1_3_11 ( .I0(ML_int_3__11_), .I1(ML_int_3__3_), .S(SH[3]), 
        .Z(ML_int_4__11_) );
  CKMUX2V2_8TH40 M1_3_10 ( .I0(ML_int_3__10_), .I1(ML_int_3__2_), .S(SH[3]), 
        .Z(ML_int_4__10_) );
  CKMUX2V2_8TH40 M1_3_9 ( .I0(ML_int_3__9_), .I1(ML_int_3__1_), .S(SH[3]), .Z(
        ML_int_4__9_) );
  CKMUX2V2_8TH40 M1_3_8 ( .I0(ML_int_3__8_), .I1(ML_int_3__0_), .S(SH[3]), .Z(
        ML_int_4__8_) );
  CKMUX2V2_8TH40 M1_3_14 ( .I0(ML_int_3__14_), .I1(ML_int_3__6_), .S(SH[3]), 
        .Z(ML_int_4__14_) );
  CKMUX2V2_8TH40 M1_3_12 ( .I0(ML_int_3__12_), .I1(ML_int_3__4_), .S(SH[3]), 
        .Z(ML_int_4__12_) );
  CKMUX2V2_8TH40 M1_2_23 ( .I0(ML_int_2__23_), .I1(ML_int_2__19_), .S(SH[2]), 
        .Z(ML_int_3__23_) );
  CKMUX2V2_8TH40 M1_2_15 ( .I0(ML_int_2__15_), .I1(ML_int_2__11_), .S(SH[2]), 
        .Z(ML_int_3__15_) );
  CKMUX2V2_8TH40 M1_2_21 ( .I0(ML_int_2__21_), .I1(ML_int_2__17_), .S(SH[2]), 
        .Z(ML_int_3__21_) );
  CKMUX2V2_8TH40 M1_2_13 ( .I0(ML_int_2__13_), .I1(ML_int_2__9_), .S(SH[2]), 
        .Z(ML_int_3__13_) );
  CKMUX2V2_8TH40 M1_2_19 ( .I0(ML_int_2__19_), .I1(ML_int_2__15_), .S(SH[2]), 
        .Z(ML_int_3__19_) );
  CKMUX2V2_8TH40 M1_2_11 ( .I0(ML_int_2__11_), .I1(ML_int_2__7_), .S(SH[2]), 
        .Z(ML_int_3__11_) );
  CKMUX2V2_8TH40 M1_2_18 ( .I0(ML_int_2__18_), .I1(ML_int_2__14_), .S(SH[2]), 
        .Z(ML_int_3__18_) );
  CKMUX2V2_8TH40 M1_2_10 ( .I0(ML_int_2__10_), .I1(ML_int_2__6_), .S(SH[2]), 
        .Z(ML_int_3__10_) );
  CKMUX2V2_8TH40 M1_2_17 ( .I0(ML_int_2__17_), .I1(ML_int_2__13_), .S(SH[2]), 
        .Z(ML_int_3__17_) );
  CKMUX2V2_8TH40 M1_2_9 ( .I0(ML_int_2__9_), .I1(ML_int_2__5_), .S(SH[2]), .Z(
        ML_int_3__9_) );
  CKMUX2V2_8TH40 M1_2_16 ( .I0(ML_int_2__16_), .I1(ML_int_2__12_), .S(SH[2]), 
        .Z(ML_int_3__16_) );
  CKMUX2V2_8TH40 M1_2_8 ( .I0(ML_int_2__8_), .I1(ML_int_2__4_), .S(SH[2]), .Z(
        ML_int_3__8_) );
  CKMUX2V2_8TH40 M1_2_22 ( .I0(ML_int_2__22_), .I1(ML_int_2__18_), .S(SH[2]), 
        .Z(ML_int_3__22_) );
  CKMUX2V2_8TH40 M1_2_14 ( .I0(ML_int_2__14_), .I1(ML_int_2__10_), .S(SH[2]), 
        .Z(ML_int_3__14_) );
  CKMUX2V2_8TH40 M1_2_20 ( .I0(ML_int_2__20_), .I1(ML_int_2__16_), .S(SH[2]), 
        .Z(ML_int_3__20_) );
  CKMUX2V2_8TH40 M1_2_12 ( .I0(ML_int_2__12_), .I1(ML_int_2__8_), .S(SH[2]), 
        .Z(ML_int_3__12_) );
  CKMUX2V2_8TH40 M1_2_7 ( .I0(ML_int_2__7_), .I1(ML_int_2__3_), .S(SH[2]), .Z(
        ML_int_3__7_) );
  CKMUX2V2_8TH40 M1_2_5 ( .I0(ML_int_2__5_), .I1(ML_int_2__1_), .S(SH[2]), .Z(
        ML_int_3__5_) );
  CKMUX2V2_8TH40 M1_2_4 ( .I0(ML_int_2__4_), .I1(ML_int_2__0_), .S(SH[2]), .Z(
        ML_int_3__4_) );
  CKMUX2V2_8TH40 M1_2_6 ( .I0(ML_int_2__6_), .I1(ML_int_2__2_), .S(SH[2]), .Z(
        ML_int_3__6_) );
  CKMUX2V2_8TH40 M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(ML_int_1__1_) );
  CKMUX2V2_8TH40 M1_0_28 ( .I0(A[28]), .I1(A[27]), .S(SH[0]), .Z(ML_int_1__28_) );
  CKMUX2V2_8TH40 M1_0_26 ( .I0(A[26]), .I1(A[25]), .S(SH[0]), .Z(ML_int_1__26_) );
  CKMUX2V2_8TH40 M1_0_24 ( .I0(A[24]), .I1(A[23]), .S(SH[0]), .Z(ML_int_1__24_) );
  CKMUX2V2_8TH40 M1_0_21 ( .I0(A[21]), .I1(A[20]), .S(SH[0]), .Z(ML_int_1__21_) );
  CKMUX2V2_8TH40 M1_0_19 ( .I0(A[19]), .I1(A[18]), .S(SH[0]), .Z(ML_int_1__19_) );
  CKMUX2V2_8TH40 M1_0_17 ( .I0(A[17]), .I1(A[16]), .S(SH[0]), .Z(ML_int_1__17_) );
  CKMUX2V2_8TH40 M1_0_15 ( .I0(A[15]), .I1(A[14]), .S(SH[0]), .Z(ML_int_1__15_) );
  CKMUX2V2_8TH40 M1_0_13 ( .I0(A[13]), .I1(A[12]), .S(SH[0]), .Z(ML_int_1__13_) );
  CKMUX2V2_8TH40 M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(ML_int_1__11_) );
  CKMUX2V2_8TH40 M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(ML_int_1__9_) );
  CKMUX2V2_8TH40 M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(ML_int_1__7_) );
  CKMUX2V2_8TH40 M1_0_29 ( .I0(A[29]), .I1(A[28]), .S(SH[0]), .Z(ML_int_1__29_) );
  CKMUX2V2_8TH40 M1_0_27 ( .I0(A[27]), .I1(A[26]), .S(SH[0]), .Z(ML_int_1__27_) );
  CKMUX2V2_8TH40 M1_0_25 ( .I0(A[25]), .I1(A[24]), .S(SH[0]), .Z(ML_int_1__25_) );
  CKMUX2V2_8TH40 M1_0_23 ( .I0(A[23]), .I1(A[22]), .S(SH[0]), .Z(ML_int_1__23_) );
  CKMUX2V2_8TH40 M1_0_22 ( .I0(A[22]), .I1(A[21]), .S(SH[0]), .Z(ML_int_1__22_) );
  CKMUX2V2_8TH40 M1_0_20 ( .I0(A[20]), .I1(A[19]), .S(SH[0]), .Z(ML_int_1__20_) );
  CKMUX2V2_8TH40 M1_0_18 ( .I0(A[18]), .I1(A[17]), .S(SH[0]), .Z(ML_int_1__18_) );
  CKMUX2V2_8TH40 M1_0_16 ( .I0(A[16]), .I1(A[15]), .S(SH[0]), .Z(ML_int_1__16_) );
  CKMUX2V2_8TH40 M1_0_14 ( .I0(A[14]), .I1(A[13]), .S(SH[0]), .Z(ML_int_1__14_) );
  CKMUX2V2_8TH40 M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(ML_int_1__12_) );
  CKMUX2V2_8TH40 M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(ML_int_1__10_)
         );
  CKMUX2V2_8TH40 M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(ML_int_1__8_) );
  CKMUX2V2_8TH40 M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(ML_int_1__5_) );
  CKMUX2V2_8TH40 M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(ML_int_1__3_) );
  CKMUX2V2_8TH40 M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(ML_int_1__2_) );
  CKMUX2V2_8TH40 M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(ML_int_1__6_) );
  CKMUX2V2_8TH40 M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(ML_int_1__4_) );
  CKMUX2V2_8TH40 M1_1_3 ( .I0(ML_int_1__3_), .I1(ML_int_1__1_), .S(SH[1]), .Z(
        ML_int_2__3_) );
  CKMUX2V2_8TH40 M1_1_2 ( .I0(ML_int_1__2_), .I1(ML_int_1__0_), .S(SH[1]), .Z(
        ML_int_2__2_) );
  CKMUX2V2_8TH40 M1_1_26 ( .I0(ML_int_1__26_), .I1(ML_int_1__24_), .S(SH[1]), 
        .Z(ML_int_2__26_) );
  CKMUX2V2_8TH40 M1_1_24 ( .I0(ML_int_1__24_), .I1(ML_int_1__22_), .S(SH[1]), 
        .Z(ML_int_2__24_) );
  CKMUX2V2_8TH40 M1_1_23 ( .I0(ML_int_1__23_), .I1(ML_int_1__21_), .S(SH[1]), 
        .Z(ML_int_2__23_) );
  CKMUX2V2_8TH40 M1_1_19 ( .I0(ML_int_1__19_), .I1(ML_int_1__17_), .S(SH[1]), 
        .Z(ML_int_2__19_) );
  CKMUX2V2_8TH40 M1_1_15 ( .I0(ML_int_1__15_), .I1(ML_int_1__13_), .S(SH[1]), 
        .Z(ML_int_2__15_) );
  CKMUX2V2_8TH40 M1_1_11 ( .I0(ML_int_1__11_), .I1(ML_int_1__9_), .S(SH[1]), 
        .Z(ML_int_2__11_) );
  CKMUX2V2_8TH40 M1_1_21 ( .I0(ML_int_1__21_), .I1(ML_int_1__19_), .S(SH[1]), 
        .Z(ML_int_2__21_) );
  CKMUX2V2_8TH40 M1_1_17 ( .I0(ML_int_1__17_), .I1(ML_int_1__15_), .S(SH[1]), 
        .Z(ML_int_2__17_) );
  CKMUX2V2_8TH40 M1_1_13 ( .I0(ML_int_1__13_), .I1(ML_int_1__11_), .S(SH[1]), 
        .Z(ML_int_2__13_) );
  CKMUX2V2_8TH40 M1_1_9 ( .I0(ML_int_1__9_), .I1(ML_int_1__7_), .S(SH[1]), .Z(
        ML_int_2__9_) );
  CKMUX2V2_8TH40 M1_1_7 ( .I0(ML_int_1__7_), .I1(ML_int_1__5_), .S(SH[1]), .Z(
        ML_int_2__7_) );
  CKMUX2V2_8TH40 M1_1_27 ( .I0(ML_int_1__27_), .I1(ML_int_1__25_), .S(SH[1]), 
        .Z(ML_int_2__27_) );
  CKMUX2V2_8TH40 M1_1_25 ( .I0(ML_int_1__25_), .I1(ML_int_1__23_), .S(SH[1]), 
        .Z(ML_int_2__25_) );
  CKMUX2V2_8TH40 M1_1_22 ( .I0(ML_int_1__22_), .I1(ML_int_1__20_), .S(SH[1]), 
        .Z(ML_int_2__22_) );
  CKMUX2V2_8TH40 M1_1_20 ( .I0(ML_int_1__20_), .I1(ML_int_1__18_), .S(SH[1]), 
        .Z(ML_int_2__20_) );
  CKMUX2V2_8TH40 M1_1_18 ( .I0(ML_int_1__18_), .I1(ML_int_1__16_), .S(SH[1]), 
        .Z(ML_int_2__18_) );
  CKMUX2V2_8TH40 M1_1_14 ( .I0(ML_int_1__14_), .I1(ML_int_1__12_), .S(SH[1]), 
        .Z(ML_int_2__14_) );
  CKMUX2V2_8TH40 M1_1_10 ( .I0(ML_int_1__10_), .I1(ML_int_1__8_), .S(SH[1]), 
        .Z(ML_int_2__10_) );
  CKMUX2V2_8TH40 M1_1_5 ( .I0(ML_int_1__5_), .I1(ML_int_1__3_), .S(SH[1]), .Z(
        ML_int_2__5_) );
  CKMUX2V2_8TH40 M1_1_16 ( .I0(ML_int_1__16_), .I1(ML_int_1__14_), .S(SH[1]), 
        .Z(ML_int_2__16_) );
  CKMUX2V2_8TH40 M1_1_12 ( .I0(ML_int_1__12_), .I1(ML_int_1__10_), .S(SH[1]), 
        .Z(ML_int_2__12_) );
  CKMUX2V2_8TH40 M1_1_8 ( .I0(ML_int_1__8_), .I1(ML_int_1__6_), .S(SH[1]), .Z(
        ML_int_2__8_) );
  CKMUX2V2_8TH40 M1_1_4 ( .I0(ML_int_1__4_), .I1(ML_int_1__2_), .S(SH[1]), .Z(
        ML_int_2__4_) );
  CKMUX2V2_8TH40 M1_1_6 ( .I0(ML_int_1__6_), .I1(ML_int_1__4_), .S(SH[1]), .Z(
        ML_int_2__6_) );
  CKMUX2V2_8TH40 M1_2_27 ( .I0(ML_int_2__27_), .I1(ML_int_2__23_), .S(SH[2]), 
        .Z(ML_int_3__27_) );
  CKMUX2V2_8TH40 M1_2_26 ( .I0(ML_int_2__26_), .I1(ML_int_2__22_), .S(SH[2]), 
        .Z(ML_int_3__26_) );
  CKMUX2V2_8TH40 M1_2_25 ( .I0(ML_int_2__25_), .I1(ML_int_2__21_), .S(SH[2]), 
        .Z(ML_int_3__25_) );
  CKMUX2V2_8TH40 M1_2_24 ( .I0(ML_int_2__24_), .I1(ML_int_2__20_), .S(SH[2]), 
        .Z(ML_int_3__24_) );
  MUX2V4_8TH40 M1_1_31 ( .I0(ML_int_1__31_), .I1(ML_int_1__29_), .S(SH[1]), 
        .Z(ML_int_2__31_) );
  MUX2V4_8TH40 M1_2_28 ( .I0(ML_int_2__28_), .I1(ML_int_2__24_), .S(SH[2]), 
        .Z(ML_int_3__28_) );
  MUX2V4_8TH40 M1_3_27 ( .I0(ML_int_3__27_), .I1(ML_int_3__19_), .S(SH[3]), 
        .Z(ML_int_4__27_) );
  MUX2V4_8TH40 M1_3_26 ( .I0(ML_int_3__26_), .I1(ML_int_3__18_), .S(SH[3]), 
        .Z(ML_int_4__26_) );
  MUX2V4_8TH40 M1_3_25 ( .I0(ML_int_3__25_), .I1(ML_int_3__17_), .S(SH[3]), 
        .Z(ML_int_4__25_) );
  MUX2V4_8TH40 M1_3_24 ( .I0(ML_int_3__24_), .I1(ML_int_3__16_), .S(SH[3]), 
        .Z(ML_int_4__24_) );
  CKMUX2V8_8TH40 M1_4_29 ( .I0(ML_int_4__29_), .I1(ML_int_4__13_), .S(SH[4]), 
        .Z(B[29]) );
  CKMUX2V8_8TH40 M1_4_27 ( .I0(ML_int_4__27_), .I1(ML_int_4__11_), .S(SH[4]), 
        .Z(B[27]) );
  CKMUX2V8_8TH40 M1_4_26 ( .I0(ML_int_4__26_), .I1(ML_int_4__10_), .S(SH[4]), 
        .Z(B[26]) );
  CKMUX2V8_8TH40 M1_4_25 ( .I0(ML_int_4__25_), .I1(ML_int_4__9_), .S(SH[4]), 
        .Z(B[25]) );
  CKMUX2V8_8TH40 M1_4_24 ( .I0(ML_int_4__24_), .I1(ML_int_4__8_), .S(SH[4]), 
        .Z(B[24]) );
  CKMUX2V8_8TH40 M1_4_31 ( .I0(ML_int_4__31_), .I1(ML_int_4__15_), .S(SH[4]), 
        .Z(B[31]) );
  CKMUX2V8_8TH40 M1_3_30 ( .I0(ML_int_3__30_), .I1(ML_int_3__22_), .S(SH[3]), 
        .Z(ML_int_4__30_) );
  CKMUX2V8_8TH40 M1_3_28 ( .I0(ML_int_3__28_), .I1(ML_int_3__20_), .S(SH[3]), 
        .Z(ML_int_4__28_) );
  CKMUX2V8_8TH40 M1_2_31 ( .I0(ML_int_2__31_), .I1(ML_int_2__27_), .S(SH[2]), 
        .Z(ML_int_3__31_) );
  CKMUX2V8_8TH40 M1_2_29 ( .I0(ML_int_2__29_), .I1(ML_int_2__25_), .S(SH[2]), 
        .Z(ML_int_3__29_) );
  CKMUX2V8_8TH40 M1_1_30 ( .I0(ML_int_1__30_), .I1(ML_int_1__28_), .S(SH[1]), 
        .Z(ML_int_2__30_) );
  MUX2NV2_8TH40 U3 ( .I0(n1), .I1(n15), .S(SH[4]), .ZN(B[20]) );
  MUX2NV2_8TH40 U4 ( .I0(n2), .I1(n13), .S(SH[4]), .ZN(B[22]) );
  MUX2NV0_8TH40 U5 ( .I0(ML_int_3__20_), .I1(ML_int_3__12_), .S(SH[3]), .ZN(n1) );
  MUX2NV0_8TH40 U6 ( .I0(ML_int_3__22_), .I1(ML_int_3__14_), .S(SH[3]), .ZN(n2) );
  INV2_8TH40 U7 ( .I(SH[3]), .ZN(n9) );
  INV2_8TH40 U8 ( .I(SH[2]), .ZN(n10) );
  INV2_8TH40 U9 ( .I(SH[1]), .ZN(n11) );
  INOR2V2_8TH40 U10 ( .A1(A[0]), .B1(SH[0]), .ZN(ML_int_1__0_) );
  MUX2NV0_8TH40 U11 ( .I0(n3), .I1(n16), .S(SH[4]), .ZN(B[19]) );
  MUX2NV0_8TH40 U12 ( .I0(ML_int_3__19_), .I1(ML_int_3__11_), .S(SH[3]), .ZN(
        n3) );
  MUX2NV0_8TH40 U13 ( .I0(n4), .I1(n12), .S(SH[4]), .ZN(B[23]) );
  MUX2NV0_8TH40 U14 ( .I0(ML_int_3__23_), .I1(ML_int_3__15_), .S(SH[3]), .ZN(
        n4) );
  MUX2NV0_8TH40 U15 ( .I0(n5), .I1(n19), .S(SH[4]), .ZN(B[16]) );
  MUX2NV0_8TH40 U16 ( .I0(ML_int_3__16_), .I1(ML_int_3__8_), .S(SH[3]), .ZN(n5) );
  MUX2NV0_8TH40 U17 ( .I0(n6), .I1(n18), .S(SH[4]), .ZN(B[17]) );
  MUX2NV0_8TH40 U18 ( .I0(ML_int_3__17_), .I1(ML_int_3__9_), .S(SH[3]), .ZN(n6) );
  MUX2NV0_8TH40 U19 ( .I0(n7), .I1(n17), .S(SH[4]), .ZN(B[18]) );
  MUX2NV0_8TH40 U20 ( .I0(ML_int_3__18_), .I1(ML_int_3__10_), .S(SH[3]), .ZN(
        n7) );
  MUX2NV0_8TH40 U21 ( .I0(n8), .I1(n14), .S(SH[4]), .ZN(B[21]) );
  MUX2NV0_8TH40 U22 ( .I0(ML_int_3__21_), .I1(ML_int_3__13_), .S(SH[3]), .ZN(
        n8) );
  INOR2V0_8TH40 U23 ( .A1(ML_int_4__9_), .B1(SH[4]), .ZN(B[9]) );
  INOR2V0_8TH40 U24 ( .A1(ML_int_4__8_), .B1(SH[4]), .ZN(B[8]) );
  NOR2V0P5_8TH40 U25 ( .A1(SH[4]), .A2(n12), .ZN(B[7]) );
  NOR2V0P5_8TH40 U26 ( .A1(SH[4]), .A2(n13), .ZN(B[6]) );
  NOR2V0P5_8TH40 U27 ( .A1(SH[4]), .A2(n14), .ZN(B[5]) );
  NOR2V0P5_8TH40 U28 ( .A1(SH[4]), .A2(n15), .ZN(B[4]) );
  NOR2V0P5_8TH40 U29 ( .A1(SH[4]), .A2(n16), .ZN(B[3]) );
  NOR2V0P5_8TH40 U30 ( .A1(SH[4]), .A2(n17), .ZN(B[2]) );
  NOR2V0P5_8TH40 U31 ( .A1(SH[4]), .A2(n18), .ZN(B[1]) );
  INOR2V0_8TH40 U32 ( .A1(ML_int_4__15_), .B1(SH[4]), .ZN(B[15]) );
  INOR2V0_8TH40 U33 ( .A1(ML_int_4__14_), .B1(SH[4]), .ZN(B[14]) );
  INOR2V0_8TH40 U34 ( .A1(ML_int_4__13_), .B1(SH[4]), .ZN(B[13]) );
  INOR2V0_8TH40 U35 ( .A1(ML_int_4__12_), .B1(SH[4]), .ZN(B[12]) );
  INOR2V0_8TH40 U36 ( .A1(ML_int_4__11_), .B1(SH[4]), .ZN(B[11]) );
  INOR2V0_8TH40 U37 ( .A1(ML_int_4__10_), .B1(SH[4]), .ZN(B[10]) );
  NOR2V0P5_8TH40 U38 ( .A1(SH[4]), .A2(n19), .ZN(B[0]) );
  CLKNAND2V1_8TH40 U39 ( .A1(ML_int_3__7_), .A2(n9), .ZN(n12) );
  CLKNAND2V1_8TH40 U40 ( .A1(ML_int_3__6_), .A2(n9), .ZN(n13) );
  CLKNAND2V1_8TH40 U41 ( .A1(ML_int_3__5_), .A2(n9), .ZN(n14) );
  CLKNAND2V1_8TH40 U42 ( .A1(ML_int_3__4_), .A2(n9), .ZN(n15) );
  CLKNAND2V1_8TH40 U43 ( .A1(ML_int_3__3_), .A2(n9), .ZN(n16) );
  CLKNAND2V1_8TH40 U44 ( .A1(ML_int_3__2_), .A2(n9), .ZN(n17) );
  CLKNAND2V1_8TH40 U45 ( .A1(ML_int_3__1_), .A2(n9), .ZN(n18) );
  CLKNAND2V1_8TH40 U46 ( .A1(ML_int_3__0_), .A2(n9), .ZN(n19) );
  AND2V0_8TH40 U47 ( .A1(ML_int_2__3_), .A2(n10), .Z(ML_int_3__3_) );
  AND2V0_8TH40 U48 ( .A1(ML_int_2__2_), .A2(n10), .Z(ML_int_3__2_) );
  AND2V0_8TH40 U49 ( .A1(ML_int_2__1_), .A2(n10), .Z(ML_int_3__1_) );
  AND2V0_8TH40 U50 ( .A1(ML_int_2__0_), .A2(n10), .Z(ML_int_3__0_) );
  AND2V0_8TH40 U51 ( .A1(ML_int_1__1_), .A2(n11), .Z(ML_int_2__1_) );
  AND2V0_8TH40 U52 ( .A1(ML_int_1__0_), .A2(n11), .Z(ML_int_2__0_) );
endmodule


module inst_execute_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126;

  NAND2V2_8TH40 U1 ( .A1(n60), .A2(n64), .ZN(n62) );
  AND2V2_8TH40 U2 ( .A1(n61), .A2(n124), .Z(n1) );
  AND2V2_8TH40 U3 ( .A1(n1), .A2(n123), .Z(n2) );
  AND2V2_8TH40 U4 ( .A1(n2), .A2(n122), .Z(n3) );
  AND2V2_8TH40 U5 ( .A1(n3), .A2(n121), .Z(n4) );
  AND2V2_8TH40 U6 ( .A1(n4), .A2(n120), .Z(n5) );
  AND2V2_8TH40 U7 ( .A1(n5), .A2(n119), .Z(n6) );
  AND2V2_8TH40 U8 ( .A1(n6), .A2(n118), .Z(n7) );
  AND2V2_8TH40 U9 ( .A1(n7), .A2(n117), .Z(n8) );
  AND2V2_8TH40 U10 ( .A1(n8), .A2(n116), .Z(n9) );
  AND2V2_8TH40 U11 ( .A1(n9), .A2(n115), .Z(n10) );
  AND2V2_8TH40 U12 ( .A1(n10), .A2(n114), .Z(n11) );
  AND2V2_8TH40 U13 ( .A1(n11), .A2(n113), .Z(n12) );
  AND2V2_8TH40 U14 ( .A1(n12), .A2(n112), .Z(n13) );
  AND2V2_8TH40 U15 ( .A1(n13), .A2(n111), .Z(n14) );
  AND2V2_8TH40 U16 ( .A1(n14), .A2(n110), .Z(n15) );
  AND2V2_8TH40 U17 ( .A1(n15), .A2(n109), .Z(n16) );
  AND2V2_8TH40 U18 ( .A1(n16), .A2(n108), .Z(n17) );
  AND2V2_8TH40 U19 ( .A1(n17), .A2(n107), .Z(n18) );
  AND2V2_8TH40 U20 ( .A1(n18), .A2(n106), .Z(n19) );
  AND2V2_8TH40 U21 ( .A1(n19), .A2(n105), .Z(n20) );
  AND2V2_8TH40 U22 ( .A1(n20), .A2(n104), .Z(n21) );
  AND2V2_8TH40 U23 ( .A1(n21), .A2(n103), .Z(n22) );
  AND2V2_8TH40 U24 ( .A1(n22), .A2(n102), .Z(n23) );
  AND2V2_8TH40 U25 ( .A1(n23), .A2(n101), .Z(n24) );
  AND2V2_8TH40 U26 ( .A1(n24), .A2(n100), .Z(n25) );
  AND2V2_8TH40 U27 ( .A1(n25), .A2(n99), .Z(n26) );
  AND2V2_8TH40 U28 ( .A1(n26), .A2(n98), .Z(n27) );
  AND2V2_8TH40 U29 ( .A1(n27), .A2(n97), .Z(n28) );
  AND2V2_8TH40 U30 ( .A1(n28), .A2(n96), .Z(n29) );
  AND2V2_8TH40 U31 ( .A1(n29), .A2(n95), .Z(n30) );
  AND2V2_8TH40 U32 ( .A1(n30), .A2(n94), .Z(n31) );
  AND2V2_8TH40 U33 ( .A1(n31), .A2(n93), .Z(n32) );
  AND2V2_8TH40 U34 ( .A1(n32), .A2(n92), .Z(n33) );
  AND2V2_8TH40 U35 ( .A1(n33), .A2(n91), .Z(n34) );
  AND2V2_8TH40 U36 ( .A1(n34), .A2(n90), .Z(n35) );
  AND2V2_8TH40 U37 ( .A1(n35), .A2(n89), .Z(n36) );
  AND2V2_8TH40 U38 ( .A1(n36), .A2(n88), .Z(n37) );
  AND2V2_8TH40 U39 ( .A1(n37), .A2(n87), .Z(n38) );
  AND2V2_8TH40 U40 ( .A1(n38), .A2(n86), .Z(n39) );
  AND2V2_8TH40 U41 ( .A1(n39), .A2(n85), .Z(n40) );
  AND2V2_8TH40 U42 ( .A1(n40), .A2(n84), .Z(n41) );
  AND2V2_8TH40 U43 ( .A1(n41), .A2(n83), .Z(n42) );
  AND2V2_8TH40 U44 ( .A1(n42), .A2(n82), .Z(n43) );
  AND2V2_8TH40 U45 ( .A1(n43), .A2(n81), .Z(n44) );
  AND2V2_8TH40 U46 ( .A1(n44), .A2(n80), .Z(n45) );
  AND2V2_8TH40 U47 ( .A1(n45), .A2(n79), .Z(n46) );
  AND2V2_8TH40 U48 ( .A1(n46), .A2(n78), .Z(n47) );
  AND2V2_8TH40 U49 ( .A1(n47), .A2(n77), .Z(n48) );
  AND2V2_8TH40 U50 ( .A1(n48), .A2(n76), .Z(n49) );
  AND2V2_8TH40 U51 ( .A1(n49), .A2(n75), .Z(n50) );
  AND2V2_8TH40 U52 ( .A1(n50), .A2(n74), .Z(n51) );
  AND2V2_8TH40 U53 ( .A1(n51), .A2(n73), .Z(n52) );
  AND2V2_8TH40 U54 ( .A1(n52), .A2(n72), .Z(n53) );
  AND2V2_8TH40 U55 ( .A1(n53), .A2(n71), .Z(n54) );
  AND2V2_8TH40 U56 ( .A1(n54), .A2(n70), .Z(n55) );
  AND2V2_8TH40 U57 ( .A1(n55), .A2(n69), .Z(n56) );
  AND2V2_8TH40 U58 ( .A1(n56), .A2(n68), .Z(n57) );
  AND2V2_8TH40 U59 ( .A1(n57), .A2(n67), .Z(n58) );
  AND2V2_8TH40 U60 ( .A1(n58), .A2(n66), .Z(n59) );
  AND2V2_8TH40 U61 ( .A1(n59), .A2(n65), .Z(n60) );
  INV2_8TH40 U62 ( .I(B[19]), .ZN(n107) );
  INV2_8TH40 U63 ( .I(B[23]), .ZN(n103) );
  INV2_8TH40 U64 ( .I(B[6]), .ZN(n120) );
  INV2_8TH40 U65 ( .I(B[8]), .ZN(n118) );
  INV2_8TH40 U66 ( .I(B[9]), .ZN(n117) );
  INV2_8TH40 U67 ( .I(B[10]), .ZN(n116) );
  INV2_8TH40 U68 ( .I(B[11]), .ZN(n115) );
  INV2_8TH40 U69 ( .I(B[13]), .ZN(n113) );
  INV2_8TH40 U70 ( .I(B[16]), .ZN(n110) );
  INV2_8TH40 U71 ( .I(B[17]), .ZN(n109) );
  INV2_8TH40 U72 ( .I(B[18]), .ZN(n108) );
  INV2_8TH40 U73 ( .I(B[21]), .ZN(n105) );
  INV2_8TH40 U74 ( .I(B[28]), .ZN(n98) );
  INV2_8TH40 U75 ( .I(B[30]), .ZN(n96) );
  INV2_8TH40 U76 ( .I(B[7]), .ZN(n119) );
  INV2_8TH40 U77 ( .I(B[15]), .ZN(n111) );
  INV2_8TH40 U78 ( .I(B[3]), .ZN(n123) );
  INV2_8TH40 U79 ( .I(B[31]), .ZN(n95) );
  INV2_8TH40 U80 ( .I(B[1]), .ZN(n125) );
  INV2_8TH40 U81 ( .I(B[2]), .ZN(n124) );
  INV2_8TH40 U82 ( .I(B[4]), .ZN(n122) );
  INV2_8TH40 U83 ( .I(B[5]), .ZN(n121) );
  INV2_8TH40 U84 ( .I(B[12]), .ZN(n114) );
  INV2_8TH40 U85 ( .I(B[14]), .ZN(n112) );
  INV2_8TH40 U86 ( .I(B[20]), .ZN(n106) );
  INV2_8TH40 U87 ( .I(B[22]), .ZN(n104) );
  INV2_8TH40 U88 ( .I(B[24]), .ZN(n102) );
  INV2_8TH40 U89 ( .I(B[25]), .ZN(n101) );
  INV2_8TH40 U90 ( .I(B[26]), .ZN(n100) );
  INV2_8TH40 U91 ( .I(B[27]), .ZN(n99) );
  INV2_8TH40 U92 ( .I(B[29]), .ZN(n97) );
  INV2_8TH40 U93 ( .I(B[32]), .ZN(n94) );
  INV2_8TH40 U94 ( .I(B[33]), .ZN(n93) );
  INV2_8TH40 U95 ( .I(B[34]), .ZN(n92) );
  INV2_8TH40 U96 ( .I(B[35]), .ZN(n91) );
  INV2_8TH40 U97 ( .I(B[36]), .ZN(n90) );
  INV2_8TH40 U98 ( .I(B[37]), .ZN(n89) );
  INV2_8TH40 U99 ( .I(B[38]), .ZN(n88) );
  INV2_8TH40 U100 ( .I(B[39]), .ZN(n87) );
  INV2_8TH40 U101 ( .I(B[40]), .ZN(n86) );
  INV2_8TH40 U102 ( .I(B[41]), .ZN(n85) );
  INV2_8TH40 U103 ( .I(B[42]), .ZN(n84) );
  INV2_8TH40 U104 ( .I(B[43]), .ZN(n83) );
  INV2_8TH40 U105 ( .I(B[44]), .ZN(n82) );
  INV2_8TH40 U106 ( .I(B[45]), .ZN(n81) );
  INV2_8TH40 U107 ( .I(B[46]), .ZN(n80) );
  INV2_8TH40 U108 ( .I(B[47]), .ZN(n79) );
  INV2_8TH40 U109 ( .I(B[48]), .ZN(n78) );
  INV2_8TH40 U110 ( .I(B[49]), .ZN(n77) );
  INV2_8TH40 U111 ( .I(B[50]), .ZN(n76) );
  INV2_8TH40 U112 ( .I(B[51]), .ZN(n75) );
  INV2_8TH40 U113 ( .I(B[52]), .ZN(n74) );
  INV2_8TH40 U114 ( .I(B[53]), .ZN(n73) );
  INV2_8TH40 U115 ( .I(B[54]), .ZN(n72) );
  INV2_8TH40 U116 ( .I(B[55]), .ZN(n71) );
  INV2_8TH40 U117 ( .I(B[56]), .ZN(n70) );
  INV2_8TH40 U118 ( .I(B[57]), .ZN(n69) );
  INV2_8TH40 U119 ( .I(B[58]), .ZN(n68) );
  INV2_8TH40 U120 ( .I(B[59]), .ZN(n67) );
  INV2_8TH40 U121 ( .I(B[60]), .ZN(n66) );
  INV2_8TH40 U122 ( .I(B[61]), .ZN(n65) );
  INV2_8TH40 U123 ( .I(B[62]), .ZN(n64) );
  INV2_8TH40 U124 ( .I(B[63]), .ZN(n63) );
  AND2V2_8TH40 U125 ( .A1(n126), .A2(n125), .Z(n61) );
  INV2_8TH40 U126 ( .I(B[0]), .ZN(n126) );
  XNOR2V2_8TH40 U127 ( .A1(n63), .A2(n62), .ZN(DIFF[63]) );
  XOR2V2_8TH40 U128 ( .A1(n60), .A2(n64), .Z(DIFF[62]) );
  XOR2V2_8TH40 U129 ( .A1(n59), .A2(n65), .Z(DIFF[61]) );
  XOR2V2_8TH40 U130 ( .A1(n58), .A2(n66), .Z(DIFF[60]) );
  XOR2V2_8TH40 U131 ( .A1(n57), .A2(n67), .Z(DIFF[59]) );
  XOR2V2_8TH40 U132 ( .A1(n56), .A2(n68), .Z(DIFF[58]) );
  XOR2V2_8TH40 U133 ( .A1(n55), .A2(n69), .Z(DIFF[57]) );
  XOR2V2_8TH40 U134 ( .A1(n54), .A2(n70), .Z(DIFF[56]) );
  XOR2V2_8TH40 U135 ( .A1(n53), .A2(n71), .Z(DIFF[55]) );
  XOR2V2_8TH40 U136 ( .A1(n52), .A2(n72), .Z(DIFF[54]) );
  XOR2V2_8TH40 U137 ( .A1(n51), .A2(n73), .Z(DIFF[53]) );
  XOR2V2_8TH40 U138 ( .A1(n50), .A2(n74), .Z(DIFF[52]) );
  XOR2V2_8TH40 U139 ( .A1(n49), .A2(n75), .Z(DIFF[51]) );
  XOR2V2_8TH40 U140 ( .A1(n48), .A2(n76), .Z(DIFF[50]) );
  XOR2V2_8TH40 U141 ( .A1(n47), .A2(n77), .Z(DIFF[49]) );
  XOR2V2_8TH40 U142 ( .A1(n46), .A2(n78), .Z(DIFF[48]) );
  XOR2V2_8TH40 U143 ( .A1(n45), .A2(n79), .Z(DIFF[47]) );
  XOR2V2_8TH40 U144 ( .A1(n44), .A2(n80), .Z(DIFF[46]) );
  XOR2V2_8TH40 U145 ( .A1(n43), .A2(n81), .Z(DIFF[45]) );
  XOR2V2_8TH40 U146 ( .A1(n42), .A2(n82), .Z(DIFF[44]) );
  XOR2V2_8TH40 U147 ( .A1(n41), .A2(n83), .Z(DIFF[43]) );
  XOR2V2_8TH40 U148 ( .A1(n40), .A2(n84), .Z(DIFF[42]) );
  XOR2V2_8TH40 U149 ( .A1(n39), .A2(n85), .Z(DIFF[41]) );
  XOR2V2_8TH40 U150 ( .A1(n38), .A2(n86), .Z(DIFF[40]) );
  XOR2V2_8TH40 U151 ( .A1(n37), .A2(n87), .Z(DIFF[39]) );
  XOR2V2_8TH40 U152 ( .A1(n36), .A2(n88), .Z(DIFF[38]) );
  XOR2V2_8TH40 U153 ( .A1(n35), .A2(n89), .Z(DIFF[37]) );
  XOR2V2_8TH40 U154 ( .A1(n34), .A2(n90), .Z(DIFF[36]) );
  XOR2V2_8TH40 U155 ( .A1(n33), .A2(n91), .Z(DIFF[35]) );
  XOR2V2_8TH40 U156 ( .A1(n32), .A2(n92), .Z(DIFF[34]) );
  XOR2V2_8TH40 U157 ( .A1(n31), .A2(n93), .Z(DIFF[33]) );
  XOR2V2_8TH40 U158 ( .A1(n30), .A2(n94), .Z(DIFF[32]) );
  XOR2V2_8TH40 U159 ( .A1(n29), .A2(n95), .Z(DIFF[31]) );
  XOR2V2_8TH40 U160 ( .A1(n28), .A2(n96), .Z(DIFF[30]) );
  XOR2V2_8TH40 U161 ( .A1(n27), .A2(n97), .Z(DIFF[29]) );
  XOR2V2_8TH40 U162 ( .A1(n26), .A2(n98), .Z(DIFF[28]) );
  XOR2V2_8TH40 U163 ( .A1(n25), .A2(n99), .Z(DIFF[27]) );
  XOR2V2_8TH40 U164 ( .A1(n24), .A2(n100), .Z(DIFF[26]) );
  XOR2V2_8TH40 U165 ( .A1(n23), .A2(n101), .Z(DIFF[25]) );
  XOR2V2_8TH40 U166 ( .A1(n22), .A2(n102), .Z(DIFF[24]) );
  XOR2V2_8TH40 U167 ( .A1(n21), .A2(n103), .Z(DIFF[23]) );
  XOR2V2_8TH40 U168 ( .A1(n20), .A2(n104), .Z(DIFF[22]) );
  XOR2V2_8TH40 U169 ( .A1(n19), .A2(n105), .Z(DIFF[21]) );
  XOR2V2_8TH40 U170 ( .A1(n18), .A2(n106), .Z(DIFF[20]) );
  XOR2V2_8TH40 U171 ( .A1(n17), .A2(n107), .Z(DIFF[19]) );
  XOR2V2_8TH40 U172 ( .A1(n16), .A2(n108), .Z(DIFF[18]) );
  XOR2V2_8TH40 U173 ( .A1(n15), .A2(n109), .Z(DIFF[17]) );
  XOR2V2_8TH40 U174 ( .A1(n14), .A2(n110), .Z(DIFF[16]) );
  XOR2V2_8TH40 U175 ( .A1(n13), .A2(n111), .Z(DIFF[15]) );
  XOR2V2_8TH40 U176 ( .A1(n12), .A2(n112), .Z(DIFF[14]) );
  XOR2V2_8TH40 U177 ( .A1(n11), .A2(n113), .Z(DIFF[13]) );
  XOR2V2_8TH40 U178 ( .A1(n10), .A2(n114), .Z(DIFF[12]) );
  XOR2V2_8TH40 U179 ( .A1(n9), .A2(n115), .Z(DIFF[11]) );
  XOR2V2_8TH40 U180 ( .A1(n8), .A2(n116), .Z(DIFF[10]) );
  XOR2V2_8TH40 U181 ( .A1(n7), .A2(n117), .Z(DIFF[9]) );
  XOR2V2_8TH40 U182 ( .A1(n6), .A2(n118), .Z(DIFF[8]) );
  XOR2V2_8TH40 U183 ( .A1(n5), .A2(n119), .Z(DIFF[7]) );
  XOR2V2_8TH40 U184 ( .A1(n4), .A2(n120), .Z(DIFF[6]) );
  XOR2V2_8TH40 U185 ( .A1(n3), .A2(n121), .Z(DIFF[5]) );
  XOR2V2_8TH40 U186 ( .A1(n2), .A2(n122), .Z(DIFF[4]) );
  XOR2V2_8TH40 U187 ( .A1(n1), .A2(n123), .Z(DIFF[3]) );
  XOR2V2_8TH40 U188 ( .A1(n61), .A2(n124), .Z(DIFF[2]) );
  XOR2V2_8TH40 U189 ( .A1(n126), .A2(n125), .Z(DIFF[1]) );
endmodule


module inst_execute_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125;
  assign DIFF[0] = B[0];

  XOR2V4_8TH40 U1 ( .A1(B[63]), .A2(n62), .Z(DIFF[63]) );
  AND2V2_8TH40 U2 ( .A1(n29), .A2(n91), .Z(n1) );
  AND2V2_8TH40 U3 ( .A1(n1), .A2(n90), .Z(n2) );
  AND2V2_8TH40 U4 ( .A1(n2), .A2(n89), .Z(n3) );
  AND2V2_8TH40 U5 ( .A1(n3), .A2(n88), .Z(n4) );
  AND2V2_8TH40 U6 ( .A1(n4), .A2(n87), .Z(n5) );
  AND2V2_8TH40 U7 ( .A1(n5), .A2(n86), .Z(n6) );
  AND2V2_8TH40 U8 ( .A1(n6), .A2(n85), .Z(n7) );
  AND2V2_8TH40 U9 ( .A1(n7), .A2(n84), .Z(n8) );
  AND2V2_8TH40 U10 ( .A1(n8), .A2(n83), .Z(n9) );
  AND2V2_8TH40 U11 ( .A1(n9), .A2(n82), .Z(n10) );
  AND2V2_8TH40 U12 ( .A1(n10), .A2(n81), .Z(n11) );
  AND2V2_8TH40 U13 ( .A1(n11), .A2(n80), .Z(n12) );
  AND2V2_8TH40 U14 ( .A1(n12), .A2(n79), .Z(n13) );
  AND2V2_8TH40 U15 ( .A1(n13), .A2(n78), .Z(n14) );
  AND2V2_8TH40 U16 ( .A1(n14), .A2(n77), .Z(n15) );
  AND2V2_8TH40 U17 ( .A1(n15), .A2(n76), .Z(n16) );
  AND2V2_8TH40 U18 ( .A1(n16), .A2(n75), .Z(n17) );
  AND2V2_8TH40 U19 ( .A1(n17), .A2(n74), .Z(n18) );
  AND2V2_8TH40 U20 ( .A1(n18), .A2(n73), .Z(n19) );
  AND2V2_8TH40 U21 ( .A1(n19), .A2(n72), .Z(n20) );
  AND2V2_8TH40 U22 ( .A1(n20), .A2(n71), .Z(n21) );
  AND2V2_8TH40 U23 ( .A1(n21), .A2(n70), .Z(n22) );
  AND2V2_8TH40 U24 ( .A1(n22), .A2(n69), .Z(n23) );
  AND2V2_8TH40 U25 ( .A1(n23), .A2(n68), .Z(n24) );
  AND2V2_8TH40 U26 ( .A1(n24), .A2(n67), .Z(n25) );
  AND2V2_8TH40 U27 ( .A1(n25), .A2(n66), .Z(n26) );
  AND2V2_8TH40 U28 ( .A1(n26), .A2(n65), .Z(n27) );
  AND2V2_8TH40 U29 ( .A1(n27), .A2(n64), .Z(n28) );
  INV2_8TH40 U30 ( .I(B[51]), .ZN(n74) );
  INV2_8TH40 U31 ( .I(B[53]), .ZN(n72) );
  INV2_8TH40 U32 ( .I(B[55]), .ZN(n70) );
  INV2_8TH40 U33 ( .I(B[57]), .ZN(n68) );
  INV2_8TH40 U34 ( .I(B[59]), .ZN(n66) );
  INV2_8TH40 U35 ( .I(B[61]), .ZN(n64) );
  NAND2V2_8TH40 U36 ( .A1(n28), .A2(n63), .ZN(n62) );
  INV2_8TH40 U37 ( .I(B[46]), .ZN(n79) );
  INV2_8TH40 U38 ( .I(B[43]), .ZN(n82) );
  INV2_8TH40 U39 ( .I(B[37]), .ZN(n88) );
  INV2_8TH40 U40 ( .I(B[40]), .ZN(n85) );
  INV2_8TH40 U41 ( .I(B[45]), .ZN(n80) );
  INV2_8TH40 U42 ( .I(B[48]), .ZN(n77) );
  INV2_8TH40 U43 ( .I(B[36]), .ZN(n89) );
  INV2_8TH40 U44 ( .I(B[39]), .ZN(n86) );
  INV2_8TH40 U45 ( .I(B[44]), .ZN(n81) );
  INV2_8TH40 U46 ( .I(B[35]), .ZN(n90) );
  INV2_8TH40 U47 ( .I(B[42]), .ZN(n83) );
  INV2_8TH40 U48 ( .I(B[47]), .ZN(n78) );
  INV2_8TH40 U49 ( .I(B[34]), .ZN(n91) );
  INV2_8TH40 U50 ( .I(B[50]), .ZN(n75) );
  INV2_8TH40 U51 ( .I(B[52]), .ZN(n73) );
  INV2_8TH40 U52 ( .I(B[54]), .ZN(n71) );
  INV2_8TH40 U53 ( .I(B[56]), .ZN(n69) );
  INV2_8TH40 U54 ( .I(B[58]), .ZN(n67) );
  INV2_8TH40 U55 ( .I(B[60]), .ZN(n65) );
  INV2_8TH40 U56 ( .I(B[41]), .ZN(n84) );
  INV2_8TH40 U57 ( .I(B[38]), .ZN(n87) );
  INV2_8TH40 U58 ( .I(B[49]), .ZN(n76) );
  AND2V2_8TH40 U59 ( .A1(n30), .A2(n92), .Z(n29) );
  INV2_8TH40 U60 ( .I(B[62]), .ZN(n63) );
  AND2V2_8TH40 U61 ( .A1(n61), .A2(n93), .Z(n30) );
  INV2_8TH40 U62 ( .I(B[33]), .ZN(n92) );
  INV2_8TH40 U63 ( .I(B[32]), .ZN(n93) );
  INV2_8TH40 U64 ( .I(B[1]), .ZN(n124) );
  AND2V2_8TH40 U65 ( .A1(n125), .A2(n124), .Z(n31) );
  AND2V2_8TH40 U66 ( .A1(n31), .A2(n123), .Z(n32) );
  AND2V2_8TH40 U67 ( .A1(n32), .A2(n122), .Z(n33) );
  AND2V2_8TH40 U68 ( .A1(n33), .A2(n121), .Z(n34) );
  AND2V2_8TH40 U69 ( .A1(n34), .A2(n120), .Z(n35) );
  AND2V2_8TH40 U70 ( .A1(n35), .A2(n119), .Z(n36) );
  AND2V2_8TH40 U71 ( .A1(n36), .A2(n118), .Z(n37) );
  AND2V2_8TH40 U72 ( .A1(n37), .A2(n117), .Z(n38) );
  AND2V2_8TH40 U73 ( .A1(n38), .A2(n116), .Z(n39) );
  AND2V2_8TH40 U74 ( .A1(n39), .A2(n115), .Z(n40) );
  AND2V2_8TH40 U75 ( .A1(n40), .A2(n114), .Z(n41) );
  AND2V2_8TH40 U76 ( .A1(n41), .A2(n113), .Z(n42) );
  AND2V2_8TH40 U77 ( .A1(n42), .A2(n112), .Z(n43) );
  AND2V2_8TH40 U78 ( .A1(n43), .A2(n111), .Z(n44) );
  AND2V2_8TH40 U79 ( .A1(n44), .A2(n110), .Z(n45) );
  AND2V2_8TH40 U80 ( .A1(n45), .A2(n109), .Z(n46) );
  AND2V2_8TH40 U81 ( .A1(n46), .A2(n108), .Z(n47) );
  AND2V2_8TH40 U82 ( .A1(n47), .A2(n107), .Z(n48) );
  AND2V2_8TH40 U83 ( .A1(n48), .A2(n106), .Z(n49) );
  AND2V2_8TH40 U84 ( .A1(n49), .A2(n105), .Z(n50) );
  AND2V2_8TH40 U85 ( .A1(n50), .A2(n104), .Z(n51) );
  AND2V2_8TH40 U86 ( .A1(n51), .A2(n103), .Z(n52) );
  AND2V2_8TH40 U87 ( .A1(n52), .A2(n102), .Z(n53) );
  AND2V2_8TH40 U88 ( .A1(n53), .A2(n101), .Z(n54) );
  AND2V2_8TH40 U89 ( .A1(n54), .A2(n100), .Z(n55) );
  AND2V2_8TH40 U90 ( .A1(n55), .A2(n99), .Z(n56) );
  AND2V2_8TH40 U91 ( .A1(n56), .A2(n98), .Z(n57) );
  AND2V2_8TH40 U92 ( .A1(n57), .A2(n97), .Z(n58) );
  AND2V2_8TH40 U93 ( .A1(n58), .A2(n96), .Z(n59) );
  AND2V2_8TH40 U94 ( .A1(n59), .A2(n95), .Z(n60) );
  AND2V2_8TH40 U95 ( .A1(n60), .A2(n94), .Z(n61) );
  INV2_8TH40 U96 ( .I(B[0]), .ZN(n125) );
  INV2_8TH40 U97 ( .I(B[2]), .ZN(n123) );
  INV2_8TH40 U98 ( .I(B[3]), .ZN(n122) );
  INV2_8TH40 U99 ( .I(B[4]), .ZN(n121) );
  INV2_8TH40 U100 ( .I(B[5]), .ZN(n120) );
  INV2_8TH40 U101 ( .I(B[6]), .ZN(n119) );
  INV2_8TH40 U102 ( .I(B[7]), .ZN(n118) );
  INV2_8TH40 U103 ( .I(B[8]), .ZN(n117) );
  INV2_8TH40 U104 ( .I(B[9]), .ZN(n116) );
  INV2_8TH40 U105 ( .I(B[10]), .ZN(n115) );
  INV2_8TH40 U106 ( .I(B[11]), .ZN(n114) );
  INV2_8TH40 U107 ( .I(B[12]), .ZN(n113) );
  INV2_8TH40 U108 ( .I(B[13]), .ZN(n112) );
  INV2_8TH40 U109 ( .I(B[14]), .ZN(n111) );
  INV2_8TH40 U110 ( .I(B[15]), .ZN(n110) );
  INV2_8TH40 U111 ( .I(B[16]), .ZN(n109) );
  INV2_8TH40 U112 ( .I(B[17]), .ZN(n108) );
  INV2_8TH40 U113 ( .I(B[18]), .ZN(n107) );
  INV2_8TH40 U114 ( .I(B[19]), .ZN(n106) );
  INV2_8TH40 U115 ( .I(B[20]), .ZN(n105) );
  INV2_8TH40 U116 ( .I(B[21]), .ZN(n104) );
  INV2_8TH40 U117 ( .I(B[22]), .ZN(n103) );
  INV2_8TH40 U118 ( .I(B[23]), .ZN(n102) );
  INV2_8TH40 U119 ( .I(B[24]), .ZN(n101) );
  INV2_8TH40 U120 ( .I(B[25]), .ZN(n100) );
  INV2_8TH40 U121 ( .I(B[26]), .ZN(n99) );
  INV2_8TH40 U122 ( .I(B[27]), .ZN(n98) );
  INV2_8TH40 U123 ( .I(B[28]), .ZN(n97) );
  INV2_8TH40 U124 ( .I(B[29]), .ZN(n96) );
  INV2_8TH40 U125 ( .I(B[30]), .ZN(n95) );
  INV2_8TH40 U126 ( .I(B[31]), .ZN(n94) );
  XOR2V2_8TH40 U127 ( .A1(n28), .A2(n63), .Z(DIFF[62]) );
  XOR2V2_8TH40 U128 ( .A1(n27), .A2(n64), .Z(DIFF[61]) );
  XOR2V2_8TH40 U129 ( .A1(n26), .A2(n65), .Z(DIFF[60]) );
  XOR2V2_8TH40 U130 ( .A1(n25), .A2(n66), .Z(DIFF[59]) );
  XOR2V2_8TH40 U131 ( .A1(n24), .A2(n67), .Z(DIFF[58]) );
  XOR2V2_8TH40 U132 ( .A1(n23), .A2(n68), .Z(DIFF[57]) );
  XOR2V2_8TH40 U133 ( .A1(n22), .A2(n69), .Z(DIFF[56]) );
  XOR2V2_8TH40 U134 ( .A1(n21), .A2(n70), .Z(DIFF[55]) );
  XOR2V2_8TH40 U135 ( .A1(n20), .A2(n71), .Z(DIFF[54]) );
  XOR2V2_8TH40 U136 ( .A1(n19), .A2(n72), .Z(DIFF[53]) );
  XOR2V2_8TH40 U137 ( .A1(n18), .A2(n73), .Z(DIFF[52]) );
  XOR2V2_8TH40 U138 ( .A1(n17), .A2(n74), .Z(DIFF[51]) );
  XOR2V2_8TH40 U139 ( .A1(n16), .A2(n75), .Z(DIFF[50]) );
  XOR2V2_8TH40 U140 ( .A1(n15), .A2(n76), .Z(DIFF[49]) );
  XOR2V2_8TH40 U141 ( .A1(n14), .A2(n77), .Z(DIFF[48]) );
  XOR2V2_8TH40 U142 ( .A1(n13), .A2(n78), .Z(DIFF[47]) );
  XOR2V2_8TH40 U143 ( .A1(n12), .A2(n79), .Z(DIFF[46]) );
  XOR2V2_8TH40 U144 ( .A1(n11), .A2(n80), .Z(DIFF[45]) );
  XOR2V2_8TH40 U145 ( .A1(n10), .A2(n81), .Z(DIFF[44]) );
  XOR2V2_8TH40 U146 ( .A1(n9), .A2(n82), .Z(DIFF[43]) );
  XOR2V2_8TH40 U147 ( .A1(n8), .A2(n83), .Z(DIFF[42]) );
  XOR2V2_8TH40 U148 ( .A1(n7), .A2(n84), .Z(DIFF[41]) );
  XOR2V2_8TH40 U149 ( .A1(n6), .A2(n85), .Z(DIFF[40]) );
  XOR2V2_8TH40 U150 ( .A1(n5), .A2(n86), .Z(DIFF[39]) );
  XOR2V2_8TH40 U151 ( .A1(n4), .A2(n87), .Z(DIFF[38]) );
  XOR2V2_8TH40 U152 ( .A1(n3), .A2(n88), .Z(DIFF[37]) );
  XOR2V2_8TH40 U153 ( .A1(n2), .A2(n89), .Z(DIFF[36]) );
  XOR2V2_8TH40 U154 ( .A1(n1), .A2(n90), .Z(DIFF[35]) );
  XOR2V2_8TH40 U155 ( .A1(n29), .A2(n91), .Z(DIFF[34]) );
  XOR2V2_8TH40 U156 ( .A1(n30), .A2(n92), .Z(DIFF[33]) );
  XOR2V2_8TH40 U157 ( .A1(n61), .A2(n93), .Z(DIFF[32]) );
  XOR2V2_8TH40 U158 ( .A1(n60), .A2(n94), .Z(DIFF[31]) );
  XOR2V2_8TH40 U159 ( .A1(n59), .A2(n95), .Z(DIFF[30]) );
  XOR2V2_8TH40 U160 ( .A1(n58), .A2(n96), .Z(DIFF[29]) );
  XOR2V2_8TH40 U161 ( .A1(n57), .A2(n97), .Z(DIFF[28]) );
  XOR2V2_8TH40 U162 ( .A1(n56), .A2(n98), .Z(DIFF[27]) );
  XOR2V2_8TH40 U163 ( .A1(n55), .A2(n99), .Z(DIFF[26]) );
  XOR2V2_8TH40 U164 ( .A1(n54), .A2(n100), .Z(DIFF[25]) );
  XOR2V2_8TH40 U165 ( .A1(n53), .A2(n101), .Z(DIFF[24]) );
  XOR2V2_8TH40 U166 ( .A1(n52), .A2(n102), .Z(DIFF[23]) );
  XOR2V2_8TH40 U167 ( .A1(n51), .A2(n103), .Z(DIFF[22]) );
  XOR2V2_8TH40 U168 ( .A1(n50), .A2(n104), .Z(DIFF[21]) );
  XOR2V2_8TH40 U169 ( .A1(n49), .A2(n105), .Z(DIFF[20]) );
  XOR2V2_8TH40 U170 ( .A1(n48), .A2(n106), .Z(DIFF[19]) );
  XOR2V2_8TH40 U171 ( .A1(n47), .A2(n107), .Z(DIFF[18]) );
  XOR2V2_8TH40 U172 ( .A1(n46), .A2(n108), .Z(DIFF[17]) );
  XOR2V2_8TH40 U173 ( .A1(n45), .A2(n109), .Z(DIFF[16]) );
  XOR2V2_8TH40 U174 ( .A1(n44), .A2(n110), .Z(DIFF[15]) );
  XOR2V2_8TH40 U175 ( .A1(n43), .A2(n111), .Z(DIFF[14]) );
  XOR2V2_8TH40 U176 ( .A1(n42), .A2(n112), .Z(DIFF[13]) );
  XOR2V2_8TH40 U177 ( .A1(n41), .A2(n113), .Z(DIFF[12]) );
  XOR2V2_8TH40 U178 ( .A1(n40), .A2(n114), .Z(DIFF[11]) );
  XOR2V2_8TH40 U179 ( .A1(n39), .A2(n115), .Z(DIFF[10]) );
  XOR2V2_8TH40 U180 ( .A1(n38), .A2(n116), .Z(DIFF[9]) );
  XOR2V2_8TH40 U181 ( .A1(n37), .A2(n117), .Z(DIFF[8]) );
  XOR2V2_8TH40 U182 ( .A1(n36), .A2(n118), .Z(DIFF[7]) );
  XOR2V2_8TH40 U183 ( .A1(n35), .A2(n119), .Z(DIFF[6]) );
  XOR2V2_8TH40 U184 ( .A1(n34), .A2(n120), .Z(DIFF[5]) );
  XOR2V2_8TH40 U185 ( .A1(n33), .A2(n121), .Z(DIFF[4]) );
  XOR2V2_8TH40 U186 ( .A1(n32), .A2(n122), .Z(DIFF[3]) );
  XOR2V2_8TH40 U187 ( .A1(n31), .A2(n123), .Z(DIFF[2]) );
  XOR2V2_8TH40 U188 ( .A1(n125), .A2(n124), .Z(DIFF[1]) );
endmodule


module inst_execute_DW01_add_0 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;
  assign SUM[30] = A[30];
  assign SUM[29] = A[29];
  assign SUM[28] = A[28];
  assign SUM[27] = A[27];
  assign SUM[26] = A[26];
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  AOAOI2111V2_8TH40 U2 ( .A1(n87), .A2(n88), .B(n89), .C(n10), .D(n9), .ZN(n81) );
  NAND4V2_8TH40 U3 ( .A1(n24), .A2(n26), .A3(n23), .A4(n143), .ZN(n92) );
  XNOR2V2_8TH40 U4 ( .A1(n73), .A2(n75), .ZN(SUM[49]) );
  XNOR2V2_8TH40 U5 ( .A1(n33), .A2(n35), .ZN(SUM[59]) );
  XNOR2V2_8TH40 U6 ( .A1(n65), .A2(n67), .ZN(SUM[51]) );
  XNOR2V2_8TH40 U7 ( .A1(n57), .A2(n59), .ZN(SUM[53]) );
  XNOR2V2_8TH40 U8 ( .A1(n49), .A2(n51), .ZN(SUM[55]) );
  XNOR2V2_8TH40 U9 ( .A1(n41), .A2(n43), .ZN(SUM[57]) );
  XOR2V2_8TH40 U10 ( .A1(n76), .A2(n79), .Z(SUM[48]) );
  AOI21V2_8TH40 U11 ( .A1(n146), .A2(n21), .B(n22), .ZN(n145) );
  AOI21V2_8TH40 U12 ( .A1(n113), .A2(n11), .B(n12), .ZN(n112) );
  XOR2V2_8TH40 U13 ( .A1(n113), .A2(n114), .Z(SUM[42]) );
  XOR2V2_8TH40 U14 ( .A1(n146), .A2(n147), .Z(SUM[34]) );
  XOR2V2_8TH40 U15 ( .A1(n131), .A2(n132), .Z(SUM[37]) );
  XOR2V2_8TH40 U16 ( .A1(n102), .A2(n117), .Z(SUM[40]) );
  XOR2V2_8TH40 U17 ( .A1(n97), .A2(n98), .Z(SUM[45]) );
  XOR2V2_8TH40 U18 ( .A1(n127), .A2(n128), .Z(SUM[39]) );
  XOR2V2_8TH40 U19 ( .A1(n68), .A2(n71), .Z(SUM[50]) );
  XOR2V2_8TH40 U20 ( .A1(n60), .A2(n63), .Z(SUM[52]) );
  XOR2V2_8TH40 U21 ( .A1(n52), .A2(n55), .Z(SUM[54]) );
  XOR2V2_8TH40 U22 ( .A1(n44), .A2(n47), .Z(SUM[56]) );
  XOR2V2_8TH40 U23 ( .A1(n36), .A2(n39), .Z(SUM[58]) );
  XOR2V2_8TH40 U24 ( .A1(n26), .A2(n151), .Z(SUM[32]) );
  XOR2V2_8TH40 U25 ( .A1(n93), .A2(n94), .Z(SUM[47]) );
  XOR2V2_8TH40 U26 ( .A1(n29), .A2(n31), .Z(SUM[60]) );
  INV2_8TH40 U27 ( .I(n90), .ZN(n9) );
  INV2_8TH40 U28 ( .I(n78), .ZN(n6) );
  INV2_8TH40 U29 ( .I(n70), .ZN(n5) );
  INV2_8TH40 U30 ( .I(n62), .ZN(n4) );
  INV2_8TH40 U31 ( .I(n54), .ZN(n3) );
  INV2_8TH40 U32 ( .I(n46), .ZN(n2) );
  INV2_8TH40 U33 ( .I(n38), .ZN(n1) );
  INV2_8TH40 U34 ( .I(n110), .ZN(n13) );
  INV2_8TH40 U35 ( .I(n120), .ZN(n17) );
  INV2_8TH40 U36 ( .I(n80), .ZN(n7) );
  INV2_8TH40 U37 ( .I(n119), .ZN(n15) );
  INV2_8TH40 U38 ( .I(n135), .ZN(n20) );
  INV2_8TH40 U39 ( .I(n139), .ZN(n21) );
  INV2_8TH40 U40 ( .I(n106), .ZN(n11) );
  INV2_8TH40 U41 ( .I(n136), .ZN(n23) );
  INV2_8TH40 U42 ( .I(n123), .ZN(n16) );
  INV2_8TH40 U43 ( .I(n150), .ZN(n24) );
  INV2_8TH40 U44 ( .I(n99), .ZN(n10) );
  INV2_8TH40 U45 ( .I(n133), .ZN(n19) );
  INV2_8TH40 U46 ( .I(n153), .ZN(n26) );
  INV2_8TH40 U47 ( .I(n137), .ZN(n25) );
  INV2_8TH40 U48 ( .I(n104), .ZN(n14) );
  INV2_8TH40 U49 ( .I(n122), .ZN(n18) );
  INV2_8TH40 U50 ( .I(n82), .ZN(n8) );
  INV2_8TH40 U51 ( .I(n140), .ZN(n22) );
  INV2_8TH40 U52 ( .I(n107), .ZN(n12) );
  INV2_8TH40 U53 ( .I(n154), .ZN(SUM[31]) );
  XNOR2V0_8TH40 U54 ( .A1(n28), .A2(B[61]), .ZN(SUM[61]) );
  OAOI211V0_8TH40 U55 ( .A1(n29), .A2(A[60]), .B(B[60]), .C(n30), .ZN(n28) );
  AND2V0_8TH40 U56 ( .A1(A[60]), .A2(n29), .Z(n30) );
  CLKXOR2V2_8TH40 U57 ( .A1(B[60]), .A2(A[60]), .Z(n31) );
  OAI21V0_8TH40 U58 ( .A1(n32), .A2(n33), .B(n34), .ZN(n29) );
  INOR2V0_8TH40 U59 ( .A1(n34), .B1(n32), .ZN(n35) );
  NOR2V0P5_8TH40 U60 ( .A1(B[59]), .A2(A[59]), .ZN(n32) );
  CLKNAND2V1_8TH40 U61 ( .A1(B[59]), .A2(A[59]), .ZN(n34) );
  AOI21V0_8TH40 U62 ( .A1(n1), .A2(n36), .B(n37), .ZN(n33) );
  NOR2V0P5_8TH40 U63 ( .A1(n37), .A2(n38), .ZN(n39) );
  NOR2V0P5_8TH40 U64 ( .A1(B[58]), .A2(A[58]), .ZN(n38) );
  AND2V0_8TH40 U65 ( .A1(B[58]), .A2(A[58]), .Z(n37) );
  OAI21V0_8TH40 U66 ( .A1(n40), .A2(n41), .B(n42), .ZN(n36) );
  INOR2V0_8TH40 U67 ( .A1(n42), .B1(n40), .ZN(n43) );
  NOR2V0P5_8TH40 U68 ( .A1(B[57]), .A2(A[57]), .ZN(n40) );
  CLKNAND2V1_8TH40 U69 ( .A1(B[57]), .A2(A[57]), .ZN(n42) );
  AOI21V0_8TH40 U70 ( .A1(n2), .A2(n44), .B(n45), .ZN(n41) );
  NOR2V0P5_8TH40 U71 ( .A1(n45), .A2(n46), .ZN(n47) );
  NOR2V0P5_8TH40 U72 ( .A1(B[56]), .A2(A[56]), .ZN(n46) );
  AND2V0_8TH40 U73 ( .A1(B[56]), .A2(A[56]), .Z(n45) );
  OAI21V0_8TH40 U74 ( .A1(n48), .A2(n49), .B(n50), .ZN(n44) );
  INOR2V0_8TH40 U75 ( .A1(n50), .B1(n48), .ZN(n51) );
  NOR2V0P5_8TH40 U76 ( .A1(B[55]), .A2(A[55]), .ZN(n48) );
  CLKNAND2V1_8TH40 U77 ( .A1(B[55]), .A2(A[55]), .ZN(n50) );
  AOI21V0_8TH40 U78 ( .A1(n3), .A2(n52), .B(n53), .ZN(n49) );
  NOR2V0P5_8TH40 U79 ( .A1(n53), .A2(n54), .ZN(n55) );
  NOR2V0P5_8TH40 U80 ( .A1(B[54]), .A2(A[54]), .ZN(n54) );
  AND2V0_8TH40 U81 ( .A1(B[54]), .A2(A[54]), .Z(n53) );
  OAI21V0_8TH40 U82 ( .A1(n56), .A2(n57), .B(n58), .ZN(n52) );
  INOR2V0_8TH40 U83 ( .A1(n58), .B1(n56), .ZN(n59) );
  NOR2V0P5_8TH40 U84 ( .A1(B[53]), .A2(A[53]), .ZN(n56) );
  CLKNAND2V1_8TH40 U85 ( .A1(B[53]), .A2(A[53]), .ZN(n58) );
  AOI21V0_8TH40 U86 ( .A1(n4), .A2(n60), .B(n61), .ZN(n57) );
  NOR2V0P5_8TH40 U87 ( .A1(n61), .A2(n62), .ZN(n63) );
  NOR2V0P5_8TH40 U88 ( .A1(B[52]), .A2(A[52]), .ZN(n62) );
  AND2V0_8TH40 U89 ( .A1(B[52]), .A2(A[52]), .Z(n61) );
  OAI21V0_8TH40 U90 ( .A1(n64), .A2(n65), .B(n66), .ZN(n60) );
  INOR2V0_8TH40 U91 ( .A1(n66), .B1(n64), .ZN(n67) );
  NOR2V0P5_8TH40 U92 ( .A1(B[51]), .A2(A[51]), .ZN(n64) );
  CLKNAND2V1_8TH40 U93 ( .A1(B[51]), .A2(A[51]), .ZN(n66) );
  AOI21V0_8TH40 U94 ( .A1(n5), .A2(n68), .B(n69), .ZN(n65) );
  NOR2V0P5_8TH40 U95 ( .A1(n69), .A2(n70), .ZN(n71) );
  NOR2V0P5_8TH40 U96 ( .A1(B[50]), .A2(A[50]), .ZN(n70) );
  AND2V0_8TH40 U97 ( .A1(B[50]), .A2(A[50]), .Z(n69) );
  OAI21V0_8TH40 U98 ( .A1(n72), .A2(n73), .B(n74), .ZN(n68) );
  INOR2V0_8TH40 U99 ( .A1(n74), .B1(n72), .ZN(n75) );
  NOR2V0P5_8TH40 U100 ( .A1(B[49]), .A2(A[49]), .ZN(n72) );
  CLKNAND2V1_8TH40 U101 ( .A1(B[49]), .A2(A[49]), .ZN(n74) );
  AOI21V0_8TH40 U102 ( .A1(n6), .A2(n76), .B(n77), .ZN(n73) );
  NOR2V0P5_8TH40 U103 ( .A1(n77), .A2(n78), .ZN(n79) );
  NOR2V0P5_8TH40 U104 ( .A1(B[48]), .A2(A[48]), .ZN(n78) );
  AND2V0_8TH40 U105 ( .A1(B[48]), .A2(A[48]), .Z(n77) );
  OAOAOAI211111V0_8TH40 U106 ( .A1(n80), .A2(n81), .B(n82), .C(n83), .D(n84), 
        .E(n85), .F(n86), .ZN(n76) );
  OAI221V0_8TH40 U107 ( .A1(n20), .A2(n91), .B1(n91), .B2(n92), .C(n15), .ZN(
        n88) );
  INOR2V0_8TH40 U108 ( .A1(n86), .B1(n85), .ZN(n94) );
  NOR2V0P5_8TH40 U109 ( .A1(B[47]), .A2(A[47]), .ZN(n85) );
  CLKNAND2V1_8TH40 U110 ( .A1(B[47]), .A2(A[47]), .ZN(n86) );
  OAI21V0_8TH40 U111 ( .A1(n83), .A2(n95), .B(n84), .ZN(n93) );
  CLKXOR2V2_8TH40 U112 ( .A1(n96), .A2(n95), .Z(SUM[46]) );
  AOI21V0_8TH40 U113 ( .A1(n7), .A2(n97), .B(n8), .ZN(n95) );
  INAND2V0_8TH40 U114 ( .A1(n83), .B1(n84), .ZN(n96) );
  CLKNAND2V1_8TH40 U115 ( .A1(B[46]), .A2(A[46]), .ZN(n84) );
  NOR2V0P5_8TH40 U116 ( .A1(B[46]), .A2(A[46]), .ZN(n83) );
  NOR2V0P5_8TH40 U117 ( .A1(n8), .A2(n80), .ZN(n98) );
  NOR2V0P5_8TH40 U118 ( .A1(B[45]), .A2(A[45]), .ZN(n80) );
  CLKNAND2V1_8TH40 U119 ( .A1(B[45]), .A2(A[45]), .ZN(n82) );
  OAI21V0_8TH40 U120 ( .A1(n99), .A2(n100), .B(n90), .ZN(n97) );
  CLKXOR2V2_8TH40 U121 ( .A1(n101), .A2(n100), .Z(SUM[44]) );
  AOI21V0_8TH40 U122 ( .A1(n102), .A2(n87), .B(n89), .ZN(n100) );
  OAOAOAI211111V0_8TH40 U123 ( .A1(n103), .A2(n104), .B(n105), .C(n106), .D(
        n107), .E(n108), .F(n109), .ZN(n89) );
  NOR4V0P5_8TH40 U124 ( .A1(n108), .A2(n106), .A3(n103), .A4(n110), .ZN(n87)
         );
  CLKNAND2V1_8TH40 U125 ( .A1(n10), .A2(n90), .ZN(n101) );
  CLKNAND2V1_8TH40 U126 ( .A1(B[44]), .A2(A[44]), .ZN(n90) );
  NOR2V0P5_8TH40 U127 ( .A1(B[44]), .A2(A[44]), .ZN(n99) );
  CLKXOR2V2_8TH40 U128 ( .A1(n111), .A2(n112), .Z(SUM[43]) );
  INAND2V0_8TH40 U129 ( .A1(n108), .B1(n109), .ZN(n111) );
  CLKNAND2V1_8TH40 U130 ( .A1(B[43]), .A2(A[43]), .ZN(n109) );
  NOR2V0P5_8TH40 U131 ( .A1(B[43]), .A2(A[43]), .ZN(n108) );
  NOR2V0P5_8TH40 U132 ( .A1(n12), .A2(n106), .ZN(n114) );
  NOR2V0P5_8TH40 U133 ( .A1(B[42]), .A2(A[42]), .ZN(n106) );
  CLKNAND2V1_8TH40 U134 ( .A1(B[42]), .A2(A[42]), .ZN(n107) );
  OAI21V0_8TH40 U135 ( .A1(n103), .A2(n115), .B(n105), .ZN(n113) );
  CLKXOR2V2_8TH40 U136 ( .A1(n116), .A2(n115), .Z(SUM[41]) );
  AOI21V0_8TH40 U137 ( .A1(n13), .A2(n102), .B(n14), .ZN(n115) );
  INAND2V0_8TH40 U138 ( .A1(n103), .B1(n105), .ZN(n116) );
  CLKNAND2V1_8TH40 U139 ( .A1(B[41]), .A2(A[41]), .ZN(n105) );
  NOR2V0P5_8TH40 U140 ( .A1(B[41]), .A2(A[41]), .ZN(n103) );
  NOR2V0P5_8TH40 U141 ( .A1(n14), .A2(n110), .ZN(n117) );
  NOR2V0P5_8TH40 U142 ( .A1(B[40]), .A2(A[40]), .ZN(n110) );
  CLKNAND2V1_8TH40 U143 ( .A1(B[40]), .A2(A[40]), .ZN(n104) );
  OAI21V0_8TH40 U144 ( .A1(n118), .A2(n91), .B(n15), .ZN(n102) );
  OAOAOAI211111V0_8TH40 U145 ( .A1(n120), .A2(n121), .B(n122), .C(n123), .D(
        n124), .E(n125), .F(n126), .ZN(n119) );
  I2NAND4V0_8TH40 U146 ( .A1(n125), .A2(n120), .B1(n16), .B2(n19), .ZN(n91) );
  INOR2V0_8TH40 U147 ( .A1(n126), .B1(n125), .ZN(n128) );
  NOR2V0P5_8TH40 U148 ( .A1(B[39]), .A2(A[39]), .ZN(n125) );
  CLKNAND2V1_8TH40 U149 ( .A1(B[39]), .A2(A[39]), .ZN(n126) );
  OAI21V0_8TH40 U150 ( .A1(n123), .A2(n129), .B(n124), .ZN(n127) );
  CLKXOR2V2_8TH40 U151 ( .A1(n130), .A2(n129), .Z(SUM[38]) );
  AOI21V0_8TH40 U152 ( .A1(n17), .A2(n131), .B(n18), .ZN(n129) );
  CLKNAND2V1_8TH40 U153 ( .A1(n16), .A2(n124), .ZN(n130) );
  CLKNAND2V1_8TH40 U154 ( .A1(B[38]), .A2(A[38]), .ZN(n124) );
  NOR2V0P5_8TH40 U155 ( .A1(B[38]), .A2(A[38]), .ZN(n123) );
  NOR2V0P5_8TH40 U156 ( .A1(n18), .A2(n120), .ZN(n132) );
  NOR2V0P5_8TH40 U157 ( .A1(B[37]), .A2(A[37]), .ZN(n120) );
  CLKNAND2V1_8TH40 U158 ( .A1(B[37]), .A2(A[37]), .ZN(n122) );
  OAI21V0_8TH40 U159 ( .A1(n133), .A2(n118), .B(n121), .ZN(n131) );
  CLKXOR2V2_8TH40 U160 ( .A1(n134), .A2(n118), .Z(SUM[36]) );
  AND2V0_8TH40 U161 ( .A1(n92), .A2(n20), .Z(n118) );
  OAOAOAI211111V0_8TH40 U162 ( .A1(n136), .A2(n137), .B(n138), .C(n139), .D(
        n140), .E(n141), .F(n142), .ZN(n135) );
  NOR2V0P5_8TH40 U163 ( .A1(n139), .A2(n141), .ZN(n143) );
  CLKNAND2V1_8TH40 U164 ( .A1(n19), .A2(n121), .ZN(n134) );
  CLKNAND2V1_8TH40 U165 ( .A1(B[36]), .A2(A[36]), .ZN(n121) );
  NOR2V0P5_8TH40 U166 ( .A1(B[36]), .A2(A[36]), .ZN(n133) );
  CLKXOR2V2_8TH40 U167 ( .A1(n144), .A2(n145), .Z(SUM[35]) );
  INAND2V0_8TH40 U168 ( .A1(n141), .B1(n142), .ZN(n144) );
  CLKNAND2V1_8TH40 U169 ( .A1(B[35]), .A2(A[35]), .ZN(n142) );
  NOR2V0P5_8TH40 U170 ( .A1(B[35]), .A2(A[35]), .ZN(n141) );
  NOR2V0P5_8TH40 U171 ( .A1(n22), .A2(n139), .ZN(n147) );
  NOR2V0P5_8TH40 U172 ( .A1(B[34]), .A2(A[34]), .ZN(n139) );
  CLKNAND2V1_8TH40 U173 ( .A1(B[34]), .A2(A[34]), .ZN(n140) );
  OAI21V0_8TH40 U174 ( .A1(n136), .A2(n148), .B(n138), .ZN(n146) );
  CLKXOR2V2_8TH40 U175 ( .A1(n149), .A2(n148), .Z(SUM[33]) );
  AOI21V0_8TH40 U176 ( .A1(n24), .A2(n26), .B(n25), .ZN(n148) );
  CLKNAND2V1_8TH40 U177 ( .A1(n23), .A2(n138), .ZN(n149) );
  CLKNAND2V1_8TH40 U178 ( .A1(B[33]), .A2(A[33]), .ZN(n138) );
  NOR2V0P5_8TH40 U179 ( .A1(B[33]), .A2(A[33]), .ZN(n136) );
  NOR2V0P5_8TH40 U180 ( .A1(n25), .A2(n150), .ZN(n151) );
  NOR2V0P5_8TH40 U181 ( .A1(B[32]), .A2(A[32]), .ZN(n150) );
  CLKNAND2V1_8TH40 U182 ( .A1(B[32]), .A2(A[32]), .ZN(n137) );
  INAND2V0_8TH40 U183 ( .A1(n152), .B1(n153), .ZN(n154) );
  CLKNAND2V1_8TH40 U184 ( .A1(B[31]), .A2(A[31]), .ZN(n153) );
  NOR2V0P5_8TH40 U185 ( .A1(B[31]), .A2(A[31]), .ZN(n152) );
endmodule


module inst_execute_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   ab_31__31_, ab_31__30_, ab_31__29_, ab_31__28_, ab_31__27_,
         ab_31__26_, ab_31__25_, ab_31__24_, ab_31__23_, ab_31__22_,
         ab_31__21_, ab_31__20_, ab_31__19_, ab_31__18_, ab_31__17_,
         ab_31__16_, ab_31__15_, ab_31__14_, ab_31__13_, ab_31__12_,
         ab_31__11_, ab_31__10_, ab_31__9_, ab_31__8_, ab_31__7_, ab_31__6_,
         ab_31__5_, ab_31__4_, ab_31__3_, ab_31__2_, ab_31__1_, ab_31__0_,
         ab_30__31_, ab_30__30_, ab_30__29_, ab_30__28_, ab_30__27_,
         ab_30__26_, ab_30__25_, ab_30__24_, ab_30__23_, ab_30__22_,
         ab_30__21_, ab_30__20_, ab_30__19_, ab_30__18_, ab_30__17_,
         ab_30__16_, ab_30__15_, ab_30__14_, ab_30__13_, ab_30__12_,
         ab_30__11_, ab_30__10_, ab_30__9_, ab_30__8_, ab_30__7_, ab_30__6_,
         ab_30__5_, ab_30__4_, ab_30__3_, ab_30__2_, ab_30__1_, ab_30__0_,
         ab_29__31_, ab_29__30_, ab_29__29_, ab_29__28_, ab_29__27_,
         ab_29__26_, ab_29__25_, ab_29__24_, ab_29__23_, ab_29__22_,
         ab_29__21_, ab_29__20_, ab_29__19_, ab_29__18_, ab_29__17_,
         ab_29__16_, ab_29__15_, ab_29__14_, ab_29__13_, ab_29__12_,
         ab_29__11_, ab_29__10_, ab_29__9_, ab_29__8_, ab_29__7_, ab_29__6_,
         ab_29__5_, ab_29__4_, ab_29__3_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__31_, ab_28__30_, ab_28__29_, ab_28__28_, ab_28__27_,
         ab_28__26_, ab_28__25_, ab_28__24_, ab_28__23_, ab_28__22_,
         ab_28__21_, ab_28__20_, ab_28__19_, ab_28__18_, ab_28__17_,
         ab_28__16_, ab_28__15_, ab_28__14_, ab_28__13_, ab_28__12_,
         ab_28__11_, ab_28__10_, ab_28__9_, ab_28__8_, ab_28__7_, ab_28__6_,
         ab_28__5_, ab_28__4_, ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_,
         ab_27__31_, ab_27__30_, ab_27__29_, ab_27__28_, ab_27__27_,
         ab_27__26_, ab_27__25_, ab_27__24_, ab_27__23_, ab_27__22_,
         ab_27__21_, ab_27__20_, ab_27__19_, ab_27__18_, ab_27__17_,
         ab_27__16_, ab_27__15_, ab_27__14_, ab_27__13_, ab_27__12_,
         ab_27__11_, ab_27__10_, ab_27__9_, ab_27__8_, ab_27__7_, ab_27__6_,
         ab_27__5_, ab_27__4_, ab_27__3_, ab_27__2_, ab_27__1_, ab_27__0_,
         ab_26__31_, ab_26__30_, ab_26__29_, ab_26__28_, ab_26__27_,
         ab_26__26_, ab_26__25_, ab_26__24_, ab_26__23_, ab_26__22_,
         ab_26__21_, ab_26__20_, ab_26__19_, ab_26__18_, ab_26__17_,
         ab_26__16_, ab_26__15_, ab_26__14_, ab_26__13_, ab_26__12_,
         ab_26__11_, ab_26__10_, ab_26__9_, ab_26__8_, ab_26__7_, ab_26__6_,
         ab_26__5_, ab_26__4_, ab_26__3_, ab_26__2_, ab_26__1_, ab_26__0_,
         ab_25__31_, ab_25__30_, ab_25__29_, ab_25__28_, ab_25__27_,
         ab_25__26_, ab_25__25_, ab_25__24_, ab_25__23_, ab_25__22_,
         ab_25__21_, ab_25__20_, ab_25__19_, ab_25__18_, ab_25__17_,
         ab_25__16_, ab_25__15_, ab_25__14_, ab_25__13_, ab_25__12_,
         ab_25__11_, ab_25__10_, ab_25__9_, ab_25__8_, ab_25__7_, ab_25__6_,
         ab_25__5_, ab_25__4_, ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_,
         ab_24__31_, ab_24__30_, ab_24__29_, ab_24__28_, ab_24__27_,
         ab_24__26_, ab_24__25_, ab_24__24_, ab_24__23_, ab_24__22_,
         ab_24__21_, ab_24__20_, ab_24__19_, ab_24__18_, ab_24__17_,
         ab_24__16_, ab_24__15_, ab_24__14_, ab_24__13_, ab_24__12_,
         ab_24__11_, ab_24__10_, ab_24__9_, ab_24__8_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__31_, ab_23__30_, ab_23__29_, ab_23__28_, ab_23__27_,
         ab_23__26_, ab_23__25_, ab_23__24_, ab_23__23_, ab_23__22_,
         ab_23__21_, ab_23__20_, ab_23__19_, ab_23__18_, ab_23__17_,
         ab_23__16_, ab_23__15_, ab_23__14_, ab_23__13_, ab_23__12_,
         ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_, ab_23__7_, ab_23__6_,
         ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_, ab_23__1_, ab_23__0_,
         ab_22__31_, ab_22__30_, ab_22__29_, ab_22__28_, ab_22__27_,
         ab_22__26_, ab_22__25_, ab_22__24_, ab_22__23_, ab_22__22_,
         ab_22__21_, ab_22__20_, ab_22__19_, ab_22__18_, ab_22__17_,
         ab_22__16_, ab_22__15_, ab_22__14_, ab_22__13_, ab_22__12_,
         ab_22__11_, ab_22__10_, ab_22__9_, ab_22__8_, ab_22__7_, ab_22__6_,
         ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_, ab_22__0_,
         ab_21__31_, ab_21__30_, ab_21__29_, ab_21__28_, ab_21__27_,
         ab_21__26_, ab_21__25_, ab_21__24_, ab_21__23_, ab_21__22_,
         ab_21__21_, ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_,
         ab_21__16_, ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_,
         ab_21__11_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__31_, ab_20__30_, ab_20__29_, ab_20__28_, ab_20__27_,
         ab_20__26_, ab_20__25_, ab_20__24_, ab_20__23_, ab_20__22_,
         ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_, ab_20__17_,
         ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_, ab_20__12_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__31_, ab_19__30_, ab_19__29_, ab_19__28_, ab_19__27_,
         ab_19__26_, ab_19__25_, ab_19__24_, ab_19__23_, ab_19__22_,
         ab_19__21_, ab_19__20_, ab_19__19_, ab_19__18_, ab_19__17_,
         ab_19__16_, ab_19__15_, ab_19__14_, ab_19__13_, ab_19__12_,
         ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_, ab_19__6_,
         ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_, ab_19__0_,
         ab_18__31_, ab_18__30_, ab_18__29_, ab_18__28_, ab_18__27_,
         ab_18__26_, ab_18__25_, ab_18__24_, ab_18__23_, ab_18__22_,
         ab_18__21_, ab_18__20_, ab_18__19_, ab_18__18_, ab_18__17_,
         ab_18__16_, ab_18__15_, ab_18__14_, ab_18__13_, ab_18__12_,
         ab_18__11_, ab_18__10_, ab_18__9_, ab_18__8_, ab_18__7_, ab_18__6_,
         ab_18__5_, ab_18__4_, ab_18__3_, ab_18__2_, ab_18__1_, ab_18__0_,
         ab_17__31_, ab_17__30_, ab_17__29_, ab_17__28_, ab_17__27_,
         ab_17__26_, ab_17__25_, ab_17__24_, ab_17__23_, ab_17__22_,
         ab_17__21_, ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_,
         ab_17__16_, ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__31_, ab_16__30_, ab_16__29_, ab_16__28_, ab_16__27_,
         ab_16__26_, ab_16__25_, ab_16__24_, ab_16__23_, ab_16__22_,
         ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_, ab_16__17_,
         ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_,
         ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_,
         ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_,
         ab_15__31_, ab_15__30_, ab_15__29_, ab_15__28_, ab_15__27_,
         ab_15__26_, ab_15__25_, ab_15__24_, ab_15__23_, ab_15__22_,
         ab_15__21_, ab_15__20_, ab_15__19_, ab_15__18_, ab_15__17_,
         ab_15__16_, ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_,
         ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_,
         ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_,
         ab_14__31_, ab_14__30_, ab_14__29_, ab_14__28_, ab_14__27_,
         ab_14__26_, ab_14__25_, ab_14__24_, ab_14__23_, ab_14__22_,
         ab_14__21_, ab_14__20_, ab_14__19_, ab_14__18_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__31_, ab_13__30_, ab_13__29_, ab_13__28_, ab_13__27_,
         ab_13__26_, ab_13__25_, ab_13__24_, ab_13__23_, ab_13__22_,
         ab_13__21_, ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_,
         ab_13__16_, ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_,
         ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_,
         ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_,
         ab_12__31_, ab_12__30_, ab_12__29_, ab_12__28_, ab_12__27_,
         ab_12__26_, ab_12__25_, ab_12__24_, ab_12__23_, ab_12__22_,
         ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_, ab_12__17_,
         ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_,
         ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_,
         ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_,
         ab_11__31_, ab_11__30_, ab_11__29_, ab_11__28_, ab_11__27_,
         ab_11__26_, ab_11__25_, ab_11__24_, ab_11__23_, ab_11__22_,
         ab_11__21_, ab_11__20_, ab_11__19_, ab_11__18_, ab_11__17_,
         ab_11__16_, ab_11__15_, ab_11__14_, ab_11__13_, ab_11__12_,
         ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__31_, ab_10__30_, ab_10__29_, ab_10__28_, ab_10__27_,
         ab_10__26_, ab_10__25_, ab_10__24_, ab_10__23_, ab_10__22_,
         ab_10__21_, ab_10__20_, ab_10__19_, ab_10__18_, ab_10__17_,
         ab_10__16_, ab_10__15_, ab_10__14_, ab_10__13_, ab_10__12_,
         ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_, ab_10__7_, ab_10__6_,
         ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_, ab_10__1_, ab_10__0_,
         ab_9__31_, ab_9__30_, ab_9__29_, ab_9__28_, ab_9__27_, ab_9__26_,
         ab_9__25_, ab_9__24_, ab_9__23_, ab_9__22_, ab_9__21_, ab_9__20_,
         ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_,
         ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_,
         ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_,
         ab_9__0_, ab_8__31_, ab_8__30_, ab_8__29_, ab_8__28_, ab_8__27_,
         ab_8__26_, ab_8__25_, ab_8__24_, ab_8__23_, ab_8__22_, ab_8__21_,
         ab_8__20_, ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_,
         ab_8__14_, ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_,
         ab_8__8_, ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_,
         ab_8__1_, ab_8__0_, ab_7__31_, ab_7__30_, ab_7__29_, ab_7__28_,
         ab_7__27_, ab_7__26_, ab_7__25_, ab_7__24_, ab_7__23_, ab_7__22_,
         ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_, ab_7__17_, ab_7__16_,
         ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_, ab_7__11_, ab_7__10_,
         ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_,
         ab_7__2_, ab_7__1_, ab_7__0_, ab_6__31_, ab_6__30_, ab_6__29_,
         ab_6__28_, ab_6__27_, ab_6__26_, ab_6__25_, ab_6__24_, ab_6__23_,
         ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_, ab_6__17_,
         ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_, ab_6__11_,
         ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_,
         ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__31_, ab_5__30_,
         ab_5__29_, ab_5__28_, ab_5__27_, ab_5__26_, ab_5__25_, ab_5__24_,
         ab_5__23_, ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_,
         ab_5__17_, ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_,
         ab_5__11_, ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_,
         ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__31_,
         ab_4__30_, ab_4__29_, ab_4__28_, ab_4__27_, ab_4__26_, ab_4__25_,
         ab_4__24_, ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_,
         ab_4__18_, ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_,
         ab_4__12_, ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_,
         ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_,
         ab_3__31_, ab_3__30_, ab_3__29_, ab_3__28_, ab_3__27_, ab_3__26_,
         ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_, ab_3__21_, ab_3__20_,
         ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_, ab_3__14_,
         ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_, ab_3__8_,
         ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_,
         ab_3__0_, ab_2__31_, ab_2__30_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__31_, ab_1__30_, ab_1__29_, ab_1__28_,
         ab_1__27_, ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_,
         ab_1__21_, ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_,
         ab_1__15_, ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_,
         ab_1__9_, ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_,
         ab_1__2_, ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_,
         ab_0__28_, ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, ab_0__1_, CARRYB_15__30_, CARRYB_15__29_,
         CARRYB_15__28_, CARRYB_15__27_, CARRYB_15__26_, CARRYB_15__25_,
         CARRYB_15__24_, CARRYB_15__23_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__30_, CARRYB_14__29_, CARRYB_14__28_,
         CARRYB_14__27_, CARRYB_14__26_, CARRYB_14__25_, CARRYB_14__24_,
         CARRYB_14__23_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__30_, CARRYB_13__29_, CARRYB_13__28_, CARRYB_13__27_,
         CARRYB_13__26_, CARRYB_13__25_, CARRYB_13__24_, CARRYB_13__23_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__30_,
         CARRYB_12__29_, CARRYB_12__28_, CARRYB_12__27_, CARRYB_12__26_,
         CARRYB_12__25_, CARRYB_12__24_, CARRYB_12__23_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__30_, CARRYB_11__29_,
         CARRYB_11__28_, CARRYB_11__27_, CARRYB_11__26_, CARRYB_11__25_,
         CARRYB_11__24_, CARRYB_11__23_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__30_, CARRYB_10__29_, CARRYB_10__28_,
         CARRYB_10__27_, CARRYB_10__26_, CARRYB_10__25_, CARRYB_10__24_,
         CARRYB_10__23_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__30_, CARRYB_9__29_, CARRYB_9__28_, CARRYB_9__27_,
         CARRYB_9__26_, CARRYB_9__25_, CARRYB_9__24_, CARRYB_9__23_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__30_, CARRYB_8__29_, CARRYB_8__28_,
         CARRYB_8__27_, CARRYB_8__26_, CARRYB_8__25_, CARRYB_8__24_,
         CARRYB_8__23_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__30_,
         CARRYB_7__29_, CARRYB_7__28_, CARRYB_7__27_, CARRYB_7__26_,
         CARRYB_7__25_, CARRYB_7__24_, CARRYB_7__23_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__30_, CARRYB_6__29_, CARRYB_6__28_, CARRYB_6__27_,
         CARRYB_6__26_, CARRYB_6__25_, CARRYB_6__24_, CARRYB_6__23_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__30_, CARRYB_5__29_, CARRYB_5__28_,
         CARRYB_5__27_, CARRYB_5__26_, CARRYB_5__25_, CARRYB_5__24_,
         CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__30_,
         CARRYB_4__29_, CARRYB_4__28_, CARRYB_4__27_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__30_, CARRYB_3__29_, CARRYB_3__28_, CARRYB_3__27_,
         CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_, CARRYB_3__23_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__30_, CARRYB_2__29_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_15__30_, SUMB_15__29_,
         SUMB_15__28_, SUMB_15__27_, SUMB_15__26_, SUMB_15__25_, SUMB_15__24_,
         SUMB_15__23_, SUMB_15__22_, SUMB_15__21_, SUMB_15__20_, SUMB_15__19_,
         SUMB_15__18_, SUMB_15__17_, SUMB_15__16_, SUMB_15__15_, SUMB_15__14_,
         SUMB_15__13_, SUMB_15__12_, SUMB_15__11_, SUMB_15__10_, SUMB_15__9_,
         SUMB_15__8_, SUMB_15__7_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__30_, SUMB_14__29_,
         SUMB_14__28_, SUMB_14__27_, SUMB_14__26_, SUMB_14__25_, SUMB_14__24_,
         SUMB_14__23_, SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_,
         SUMB_14__18_, SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_,
         SUMB_14__13_, SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_,
         SUMB_14__8_, SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_,
         SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__30_, SUMB_13__29_,
         SUMB_13__28_, SUMB_13__27_, SUMB_13__26_, SUMB_13__25_, SUMB_13__24_,
         SUMB_13__23_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_, SUMB_13__19_,
         SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_, SUMB_13__14_,
         SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_, SUMB_13__9_,
         SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_,
         SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__30_, SUMB_12__29_,
         SUMB_12__28_, SUMB_12__27_, SUMB_12__26_, SUMB_12__25_, SUMB_12__24_,
         SUMB_12__23_, SUMB_12__22_, SUMB_12__21_, SUMB_12__20_, SUMB_12__19_,
         SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_, SUMB_12__14_,
         SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_, SUMB_12__9_,
         SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__30_, SUMB_11__29_,
         SUMB_11__28_, SUMB_11__27_, SUMB_11__26_, SUMB_11__25_, SUMB_11__24_,
         SUMB_11__23_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__30_, SUMB_10__29_,
         SUMB_10__28_, SUMB_10__27_, SUMB_10__26_, SUMB_10__25_, SUMB_10__24_,
         SUMB_10__23_, SUMB_10__22_, SUMB_10__21_, SUMB_10__20_, SUMB_10__19_,
         SUMB_10__18_, SUMB_10__17_, SUMB_10__16_, SUMB_10__15_, SUMB_10__14_,
         SUMB_10__13_, SUMB_10__12_, SUMB_10__11_, SUMB_10__10_, SUMB_10__9_,
         SUMB_10__8_, SUMB_10__7_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__30_, SUMB_9__29_,
         SUMB_9__28_, SUMB_9__27_, SUMB_9__26_, SUMB_9__25_, SUMB_9__24_,
         SUMB_9__23_, SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_,
         SUMB_9__18_, SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_,
         SUMB_9__13_, SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_,
         SUMB_9__8_, SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_,
         SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__30_, SUMB_8__29_,
         SUMB_8__28_, SUMB_8__27_, SUMB_8__26_, SUMB_8__25_, SUMB_8__24_,
         SUMB_8__23_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_, SUMB_8__19_,
         SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_, SUMB_8__14_,
         SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_, SUMB_8__9_,
         SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_,
         SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__30_, SUMB_7__29_,
         SUMB_7__28_, SUMB_7__27_, SUMB_7__26_, SUMB_7__25_, SUMB_7__24_,
         SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_, SUMB_7__19_,
         SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_, SUMB_7__14_,
         SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_, SUMB_7__9_,
         SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__30_, SUMB_6__29_,
         SUMB_6__28_, SUMB_6__27_, SUMB_6__26_, SUMB_6__25_, SUMB_6__24_,
         SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__30_, SUMB_5__29_,
         SUMB_5__28_, SUMB_5__27_, SUMB_5__26_, SUMB_5__25_, SUMB_5__24_,
         SUMB_5__23_, SUMB_5__22_, SUMB_5__21_, SUMB_5__20_, SUMB_5__19_,
         SUMB_5__18_, SUMB_5__17_, SUMB_5__16_, SUMB_5__15_, SUMB_5__14_,
         SUMB_5__13_, SUMB_5__12_, SUMB_5__11_, SUMB_5__10_, SUMB_5__9_,
         SUMB_5__8_, SUMB_5__7_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__30_, SUMB_4__29_,
         SUMB_4__28_, SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_,
         SUMB_4__23_, SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_,
         SUMB_4__18_, SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_,
         SUMB_4__13_, SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_,
         SUMB_4__8_, SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_,
         SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__30_, SUMB_3__29_,
         SUMB_3__28_, SUMB_3__27_, SUMB_3__26_, SUMB_3__25_, SUMB_3__24_,
         SUMB_3__23_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_, SUMB_3__19_,
         SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_, SUMB_3__14_,
         SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_, SUMB_3__9_,
         SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_,
         SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__30_, SUMB_2__29_,
         SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_, SUMB_2__24_,
         SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_, SUMB_2__19_,
         SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_, SUMB_2__14_,
         SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_, SUMB_2__9_,
         SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__30_, SUMB_1__29_,
         SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_, SUMB_1__24_,
         SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_31__30_, CARRYB_31__29_,
         CARRYB_31__28_, CARRYB_31__27_, CARRYB_31__26_, CARRYB_31__25_,
         CARRYB_31__24_, CARRYB_31__23_, CARRYB_31__22_, CARRYB_31__21_,
         CARRYB_31__20_, CARRYB_31__19_, CARRYB_31__18_, CARRYB_31__17_,
         CARRYB_31__16_, CARRYB_31__15_, CARRYB_31__14_, CARRYB_31__13_,
         CARRYB_31__12_, CARRYB_31__11_, CARRYB_31__10_, CARRYB_31__9_,
         CARRYB_31__8_, CARRYB_31__7_, CARRYB_31__6_, CARRYB_31__5_,
         CARRYB_31__4_, CARRYB_31__3_, CARRYB_31__2_, CARRYB_31__1_,
         CARRYB_31__0_, CARRYB_30__30_, CARRYB_30__29_, CARRYB_30__28_,
         CARRYB_30__27_, CARRYB_30__26_, CARRYB_30__25_, CARRYB_30__24_,
         CARRYB_30__23_, CARRYB_30__22_, CARRYB_30__21_, CARRYB_30__20_,
         CARRYB_30__19_, CARRYB_30__18_, CARRYB_30__17_, CARRYB_30__16_,
         CARRYB_30__15_, CARRYB_30__14_, CARRYB_30__13_, CARRYB_30__12_,
         CARRYB_30__11_, CARRYB_30__10_, CARRYB_30__9_, CARRYB_30__8_,
         CARRYB_30__7_, CARRYB_30__6_, CARRYB_30__5_, CARRYB_30__4_,
         CARRYB_30__3_, CARRYB_30__2_, CARRYB_30__1_, CARRYB_30__0_,
         CARRYB_29__30_, CARRYB_29__29_, CARRYB_29__28_, CARRYB_29__27_,
         CARRYB_29__26_, CARRYB_29__25_, CARRYB_29__24_, CARRYB_29__23_,
         CARRYB_29__22_, CARRYB_29__21_, CARRYB_29__20_, CARRYB_29__19_,
         CARRYB_29__18_, CARRYB_29__17_, CARRYB_29__16_, CARRYB_29__15_,
         CARRYB_29__14_, CARRYB_29__13_, CARRYB_29__12_, CARRYB_29__11_,
         CARRYB_29__10_, CARRYB_29__9_, CARRYB_29__8_, CARRYB_29__7_,
         CARRYB_29__6_, CARRYB_29__5_, CARRYB_29__4_, CARRYB_29__3_,
         CARRYB_29__2_, CARRYB_29__1_, CARRYB_29__0_, CARRYB_28__30_,
         CARRYB_28__29_, CARRYB_28__28_, CARRYB_28__27_, CARRYB_28__26_,
         CARRYB_28__25_, CARRYB_28__24_, CARRYB_28__23_, CARRYB_28__22_,
         CARRYB_28__21_, CARRYB_28__20_, CARRYB_28__19_, CARRYB_28__18_,
         CARRYB_28__17_, CARRYB_28__16_, CARRYB_28__15_, CARRYB_28__14_,
         CARRYB_28__13_, CARRYB_28__12_, CARRYB_28__11_, CARRYB_28__10_,
         CARRYB_28__9_, CARRYB_28__8_, CARRYB_28__7_, CARRYB_28__6_,
         CARRYB_28__5_, CARRYB_28__4_, CARRYB_28__3_, CARRYB_28__2_,
         CARRYB_28__1_, CARRYB_28__0_, CARRYB_27__30_, CARRYB_27__29_,
         CARRYB_27__28_, CARRYB_27__27_, CARRYB_27__26_, CARRYB_27__25_,
         CARRYB_27__24_, CARRYB_27__23_, CARRYB_27__22_, CARRYB_27__21_,
         CARRYB_27__20_, CARRYB_27__19_, CARRYB_27__18_, CARRYB_27__17_,
         CARRYB_27__16_, CARRYB_27__15_, CARRYB_27__14_, CARRYB_27__13_,
         CARRYB_27__12_, CARRYB_27__11_, CARRYB_27__10_, CARRYB_27__9_,
         CARRYB_27__8_, CARRYB_27__7_, CARRYB_27__6_, CARRYB_27__5_,
         CARRYB_27__4_, CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_,
         CARRYB_27__0_, CARRYB_26__30_, CARRYB_26__29_, CARRYB_26__28_,
         CARRYB_26__27_, CARRYB_26__26_, CARRYB_26__25_, CARRYB_26__24_,
         CARRYB_26__23_, CARRYB_26__22_, CARRYB_26__21_, CARRYB_26__20_,
         CARRYB_26__19_, CARRYB_26__18_, CARRYB_26__17_, CARRYB_26__16_,
         CARRYB_26__15_, CARRYB_26__14_, CARRYB_26__13_, CARRYB_26__12_,
         CARRYB_26__11_, CARRYB_26__10_, CARRYB_26__9_, CARRYB_26__8_,
         CARRYB_26__7_, CARRYB_26__6_, CARRYB_26__5_, CARRYB_26__4_,
         CARRYB_26__3_, CARRYB_26__2_, CARRYB_26__1_, CARRYB_26__0_,
         CARRYB_25__30_, CARRYB_25__29_, CARRYB_25__28_, CARRYB_25__27_,
         CARRYB_25__26_, CARRYB_25__25_, CARRYB_25__24_, CARRYB_25__23_,
         CARRYB_25__22_, CARRYB_25__21_, CARRYB_25__20_, CARRYB_25__19_,
         CARRYB_25__18_, CARRYB_25__17_, CARRYB_25__16_, CARRYB_25__15_,
         CARRYB_25__14_, CARRYB_25__13_, CARRYB_25__12_, CARRYB_25__11_,
         CARRYB_25__10_, CARRYB_25__9_, CARRYB_25__8_, CARRYB_25__7_,
         CARRYB_25__6_, CARRYB_25__5_, CARRYB_25__4_, CARRYB_25__3_,
         CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_, CARRYB_24__30_,
         CARRYB_24__29_, CARRYB_24__28_, CARRYB_24__27_, CARRYB_24__26_,
         CARRYB_24__25_, CARRYB_24__24_, CARRYB_24__23_, CARRYB_24__22_,
         CARRYB_24__21_, CARRYB_24__20_, CARRYB_24__19_, CARRYB_24__18_,
         CARRYB_24__17_, CARRYB_24__16_, CARRYB_24__15_, CARRYB_24__14_,
         CARRYB_24__13_, CARRYB_24__12_, CARRYB_24__11_, CARRYB_24__10_,
         CARRYB_24__9_, CARRYB_24__8_, CARRYB_24__7_, CARRYB_24__6_,
         CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_, CARRYB_24__2_,
         CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__30_, CARRYB_23__29_,
         CARRYB_23__28_, CARRYB_23__27_, CARRYB_23__26_, CARRYB_23__25_,
         CARRYB_23__24_, CARRYB_23__23_, CARRYB_23__22_, CARRYB_23__21_,
         CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_,
         CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_,
         CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_,
         CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__30_, CARRYB_22__29_, CARRYB_22__28_,
         CARRYB_22__27_, CARRYB_22__26_, CARRYB_22__25_, CARRYB_22__24_,
         CARRYB_22__23_, CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_,
         CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_,
         CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_,
         CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__30_, CARRYB_21__29_, CARRYB_21__28_, CARRYB_21__27_,
         CARRYB_21__26_, CARRYB_21__25_, CARRYB_21__24_, CARRYB_21__23_,
         CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_,
         CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_,
         CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_,
         CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__30_,
         CARRYB_20__29_, CARRYB_20__28_, CARRYB_20__27_, CARRYB_20__26_,
         CARRYB_20__25_, CARRYB_20__24_, CARRYB_20__23_, CARRYB_20__22_,
         CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_,
         CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_,
         CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__30_, CARRYB_19__29_,
         CARRYB_19__28_, CARRYB_19__27_, CARRYB_19__26_, CARRYB_19__25_,
         CARRYB_19__24_, CARRYB_19__23_, CARRYB_19__22_, CARRYB_19__21_,
         CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_,
         CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_,
         CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__30_, CARRYB_18__29_, CARRYB_18__28_,
         CARRYB_18__27_, CARRYB_18__26_, CARRYB_18__25_, CARRYB_18__24_,
         CARRYB_18__23_, CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_,
         CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_,
         CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__30_, CARRYB_17__29_, CARRYB_17__28_, CARRYB_17__27_,
         CARRYB_17__26_, CARRYB_17__25_, CARRYB_17__24_, CARRYB_17__23_,
         CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_,
         CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_,
         CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__30_,
         CARRYB_16__29_, CARRYB_16__28_, CARRYB_16__27_, CARRYB_16__26_,
         CARRYB_16__25_, CARRYB_16__24_, CARRYB_16__23_, CARRYB_16__22_,
         CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_,
         CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, SUMB_31__30_, SUMB_31__29_,
         SUMB_31__28_, SUMB_31__27_, SUMB_31__26_, SUMB_31__25_, SUMB_31__24_,
         SUMB_31__23_, SUMB_31__22_, SUMB_31__21_, SUMB_31__20_, SUMB_31__19_,
         SUMB_31__18_, SUMB_31__17_, SUMB_31__16_, SUMB_31__15_, SUMB_31__14_,
         SUMB_31__13_, SUMB_31__12_, SUMB_31__11_, SUMB_31__10_, SUMB_31__9_,
         SUMB_31__8_, SUMB_31__7_, SUMB_31__6_, SUMB_31__5_, SUMB_31__4_,
         SUMB_31__3_, SUMB_31__2_, SUMB_31__1_, SUMB_31__0_, SUMB_30__30_,
         SUMB_30__29_, SUMB_30__28_, SUMB_30__27_, SUMB_30__26_, SUMB_30__25_,
         SUMB_30__24_, SUMB_30__23_, SUMB_30__22_, SUMB_30__21_, SUMB_30__20_,
         SUMB_30__19_, SUMB_30__18_, SUMB_30__17_, SUMB_30__16_, SUMB_30__15_,
         SUMB_30__14_, SUMB_30__13_, SUMB_30__12_, SUMB_30__11_, SUMB_30__10_,
         SUMB_30__9_, SUMB_30__8_, SUMB_30__7_, SUMB_30__6_, SUMB_30__5_,
         SUMB_30__4_, SUMB_30__3_, SUMB_30__2_, SUMB_30__1_, SUMB_29__30_,
         SUMB_29__29_, SUMB_29__28_, SUMB_29__27_, SUMB_29__26_, SUMB_29__25_,
         SUMB_29__24_, SUMB_29__23_, SUMB_29__22_, SUMB_29__21_, SUMB_29__20_,
         SUMB_29__19_, SUMB_29__18_, SUMB_29__17_, SUMB_29__16_, SUMB_29__15_,
         SUMB_29__14_, SUMB_29__13_, SUMB_29__12_, SUMB_29__11_, SUMB_29__10_,
         SUMB_29__9_, SUMB_29__8_, SUMB_29__7_, SUMB_29__6_, SUMB_29__5_,
         SUMB_29__4_, SUMB_29__3_, SUMB_29__2_, SUMB_29__1_, SUMB_28__30_,
         SUMB_28__29_, SUMB_28__28_, SUMB_28__27_, SUMB_28__26_, SUMB_28__25_,
         SUMB_28__24_, SUMB_28__23_, SUMB_28__22_, SUMB_28__21_, SUMB_28__20_,
         SUMB_28__19_, SUMB_28__18_, SUMB_28__17_, SUMB_28__16_, SUMB_28__15_,
         SUMB_28__14_, SUMB_28__13_, SUMB_28__12_, SUMB_28__11_, SUMB_28__10_,
         SUMB_28__9_, SUMB_28__8_, SUMB_28__7_, SUMB_28__6_, SUMB_28__5_,
         SUMB_28__4_, SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__30_,
         SUMB_27__29_, SUMB_27__28_, SUMB_27__27_, SUMB_27__26_, SUMB_27__25_,
         SUMB_27__24_, SUMB_27__23_, SUMB_27__22_, SUMB_27__21_, SUMB_27__20_,
         SUMB_27__19_, SUMB_27__18_, SUMB_27__17_, SUMB_27__16_, SUMB_27__15_,
         SUMB_27__14_, SUMB_27__13_, SUMB_27__12_, SUMB_27__11_, SUMB_27__10_,
         SUMB_27__9_, SUMB_27__8_, SUMB_27__7_, SUMB_27__6_, SUMB_27__5_,
         SUMB_27__4_, SUMB_27__3_, SUMB_27__2_, SUMB_27__1_, SUMB_26__30_,
         SUMB_26__29_, SUMB_26__28_, SUMB_26__27_, SUMB_26__26_, SUMB_26__25_,
         SUMB_26__24_, SUMB_26__23_, SUMB_26__22_, SUMB_26__21_, SUMB_26__20_,
         SUMB_26__19_, SUMB_26__18_, SUMB_26__17_, SUMB_26__16_, SUMB_26__15_,
         SUMB_26__14_, SUMB_26__13_, SUMB_26__12_, SUMB_26__11_, SUMB_26__10_,
         SUMB_26__9_, SUMB_26__8_, SUMB_26__7_, SUMB_26__6_, SUMB_26__5_,
         SUMB_26__4_, SUMB_26__3_, SUMB_26__2_, SUMB_26__1_, SUMB_25__30_,
         SUMB_25__29_, SUMB_25__28_, SUMB_25__27_, SUMB_25__26_, SUMB_25__25_,
         SUMB_25__24_, SUMB_25__23_, SUMB_25__22_, SUMB_25__21_, SUMB_25__20_,
         SUMB_25__19_, SUMB_25__18_, SUMB_25__17_, SUMB_25__16_, SUMB_25__15_,
         SUMB_25__14_, SUMB_25__13_, SUMB_25__12_, SUMB_25__11_, SUMB_25__10_,
         SUMB_25__9_, SUMB_25__8_, SUMB_25__7_, SUMB_25__6_, SUMB_25__5_,
         SUMB_25__4_, SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__30_,
         SUMB_24__29_, SUMB_24__28_, SUMB_24__27_, SUMB_24__26_, SUMB_24__25_,
         SUMB_24__24_, SUMB_24__23_, SUMB_24__22_, SUMB_24__21_, SUMB_24__20_,
         SUMB_24__19_, SUMB_24__18_, SUMB_24__17_, SUMB_24__16_, SUMB_24__15_,
         SUMB_24__14_, SUMB_24__13_, SUMB_24__12_, SUMB_24__11_, SUMB_24__10_,
         SUMB_24__9_, SUMB_24__8_, SUMB_24__7_, SUMB_24__6_, SUMB_24__5_,
         SUMB_24__4_, SUMB_24__3_, SUMB_24__2_, SUMB_24__1_, SUMB_23__30_,
         SUMB_23__29_, SUMB_23__28_, SUMB_23__27_, SUMB_23__26_, SUMB_23__25_,
         SUMB_23__24_, SUMB_23__23_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_,
         SUMB_23__19_, SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_,
         SUMB_23__14_, SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_,
         SUMB_23__9_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__30_,
         SUMB_22__29_, SUMB_22__28_, SUMB_22__27_, SUMB_22__26_, SUMB_22__25_,
         SUMB_22__24_, SUMB_22__23_, SUMB_22__22_, SUMB_22__21_, SUMB_22__20_,
         SUMB_22__19_, SUMB_22__18_, SUMB_22__17_, SUMB_22__16_, SUMB_22__15_,
         SUMB_22__14_, SUMB_22__13_, SUMB_22__12_, SUMB_22__11_, SUMB_22__10_,
         SUMB_22__9_, SUMB_22__8_, SUMB_22__7_, SUMB_22__6_, SUMB_22__5_,
         SUMB_22__4_, SUMB_22__3_, SUMB_22__2_, SUMB_22__1_, SUMB_21__30_,
         SUMB_21__29_, SUMB_21__28_, SUMB_21__27_, SUMB_21__26_, SUMB_21__25_,
         SUMB_21__24_, SUMB_21__23_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_,
         SUMB_21__19_, SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_,
         SUMB_21__14_, SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_,
         SUMB_21__9_, SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_,
         SUMB_21__4_, SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__30_,
         SUMB_20__29_, SUMB_20__28_, SUMB_20__27_, SUMB_20__26_, SUMB_20__25_,
         SUMB_20__24_, SUMB_20__23_, SUMB_20__22_, SUMB_20__21_, SUMB_20__20_,
         SUMB_20__19_, SUMB_20__18_, SUMB_20__17_, SUMB_20__16_, SUMB_20__15_,
         SUMB_20__14_, SUMB_20__13_, SUMB_20__12_, SUMB_20__11_, SUMB_20__10_,
         SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_,
         SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__30_,
         SUMB_19__29_, SUMB_19__28_, SUMB_19__27_, SUMB_19__26_, SUMB_19__25_,
         SUMB_19__24_, SUMB_19__23_, SUMB_19__22_, SUMB_19__21_, SUMB_19__20_,
         SUMB_19__19_, SUMB_19__18_, SUMB_19__17_, SUMB_19__16_, SUMB_19__15_,
         SUMB_19__14_, SUMB_19__13_, SUMB_19__12_, SUMB_19__11_, SUMB_19__10_,
         SUMB_19__9_, SUMB_19__8_, SUMB_19__7_, SUMB_19__6_, SUMB_19__5_,
         SUMB_19__4_, SUMB_19__3_, SUMB_19__2_, SUMB_19__1_, SUMB_18__30_,
         SUMB_18__29_, SUMB_18__28_, SUMB_18__27_, SUMB_18__26_, SUMB_18__25_,
         SUMB_18__24_, SUMB_18__23_, SUMB_18__22_, SUMB_18__21_, SUMB_18__20_,
         SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_, SUMB_18__15_,
         SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__30_,
         SUMB_17__29_, SUMB_17__28_, SUMB_17__27_, SUMB_17__26_, SUMB_17__25_,
         SUMB_17__24_, SUMB_17__23_, SUMB_17__22_, SUMB_17__21_, SUMB_17__20_,
         SUMB_17__19_, SUMB_17__18_, SUMB_17__17_, SUMB_17__16_, SUMB_17__15_,
         SUMB_17__14_, SUMB_17__13_, SUMB_17__12_, SUMB_17__11_, SUMB_17__10_,
         SUMB_17__9_, SUMB_17__8_, SUMB_17__7_, SUMB_17__6_, SUMB_17__5_,
         SUMB_17__4_, SUMB_17__3_, SUMB_17__2_, SUMB_17__1_, SUMB_16__30_,
         SUMB_16__29_, SUMB_16__28_, SUMB_16__27_, SUMB_16__26_, SUMB_16__25_,
         SUMB_16__24_, SUMB_16__23_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_,
         SUMB_16__19_, SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_,
         SUMB_16__14_, SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_,
         SUMB_16__9_, SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_,
         SUMB_16__4_, SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, A1_60_, A1_59_,
         A1_58_, A1_57_, A1_56_, A1_55_, A1_54_, A1_53_, A1_52_, A1_51_,
         A1_50_, A1_49_, A1_48_, A1_47_, A1_46_, A1_45_, A1_44_, A1_43_,
         A1_42_, A1_41_, A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_,
         A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, A1_28_, A1_27_, A1_26_,
         A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127;

  AD1V2C_8TH40 S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .CO(
        CARRYB_31__0_), .S(SUMB_31__0_) );
  AD1V2C_8TH40 S4_1 ( .A(ab_31__1_), .B(CARRYB_30__1_), .CI(SUMB_30__2_), .CO(
        CARRYB_31__1_), .S(SUMB_31__1_) );
  AD1V2C_8TH40 S4_2 ( .A(ab_31__2_), .B(CARRYB_30__2_), .CI(SUMB_30__3_), .CO(
        CARRYB_31__2_), .S(SUMB_31__2_) );
  AD1V2C_8TH40 S4_3 ( .A(ab_31__3_), .B(CARRYB_30__3_), .CI(SUMB_30__4_), .CO(
        CARRYB_31__3_), .S(SUMB_31__3_) );
  AD1V2C_8TH40 S4_4 ( .A(ab_31__4_), .B(CARRYB_30__4_), .CI(SUMB_30__5_), .CO(
        CARRYB_31__4_), .S(SUMB_31__4_) );
  AD1V2C_8TH40 S4_5 ( .A(ab_31__5_), .B(CARRYB_30__5_), .CI(SUMB_30__6_), .CO(
        CARRYB_31__5_), .S(SUMB_31__5_) );
  AD1V2C_8TH40 S4_6 ( .A(ab_31__6_), .B(CARRYB_30__6_), .CI(SUMB_30__7_), .CO(
        CARRYB_31__6_), .S(SUMB_31__6_) );
  AD1V2C_8TH40 S4_7 ( .A(ab_31__7_), .B(CARRYB_30__7_), .CI(SUMB_30__8_), .CO(
        CARRYB_31__7_), .S(SUMB_31__7_) );
  AD1V2C_8TH40 S4_8 ( .A(ab_31__8_), .B(CARRYB_30__8_), .CI(SUMB_30__9_), .CO(
        CARRYB_31__8_), .S(SUMB_31__8_) );
  AD1V2C_8TH40 S4_9 ( .A(ab_31__9_), .B(CARRYB_30__9_), .CI(SUMB_30__10_), 
        .CO(CARRYB_31__9_), .S(SUMB_31__9_) );
  AD1V2C_8TH40 S4_10 ( .A(ab_31__10_), .B(CARRYB_30__10_), .CI(SUMB_30__11_), 
        .CO(CARRYB_31__10_), .S(SUMB_31__10_) );
  AD1V2C_8TH40 S4_11 ( .A(ab_31__11_), .B(CARRYB_30__11_), .CI(SUMB_30__12_), 
        .CO(CARRYB_31__11_), .S(SUMB_31__11_) );
  AD1V2C_8TH40 S4_12 ( .A(ab_31__12_), .B(CARRYB_30__12_), .CI(SUMB_30__13_), 
        .CO(CARRYB_31__12_), .S(SUMB_31__12_) );
  AD1V2C_8TH40 S4_13 ( .A(ab_31__13_), .B(CARRYB_30__13_), .CI(SUMB_30__14_), 
        .CO(CARRYB_31__13_), .S(SUMB_31__13_) );
  AD1V2C_8TH40 S4_14 ( .A(ab_31__14_), .B(CARRYB_30__14_), .CI(SUMB_30__15_), 
        .CO(CARRYB_31__14_), .S(SUMB_31__14_) );
  AD1V2C_8TH40 S4_15 ( .A(ab_31__15_), .B(CARRYB_30__15_), .CI(SUMB_30__16_), 
        .CO(CARRYB_31__15_), .S(SUMB_31__15_) );
  AD1V2C_8TH40 S4_16 ( .A(ab_31__16_), .B(CARRYB_30__16_), .CI(SUMB_30__17_), 
        .CO(CARRYB_31__16_), .S(SUMB_31__16_) );
  AD1V2C_8TH40 S4_17 ( .A(ab_31__17_), .B(CARRYB_30__17_), .CI(SUMB_30__18_), 
        .CO(CARRYB_31__17_), .S(SUMB_31__17_) );
  AD1V2C_8TH40 S4_18 ( .A(ab_31__18_), .B(CARRYB_30__18_), .CI(SUMB_30__19_), 
        .CO(CARRYB_31__18_), .S(SUMB_31__18_) );
  AD1V2C_8TH40 S4_19 ( .A(ab_31__19_), .B(CARRYB_30__19_), .CI(SUMB_30__20_), 
        .CO(CARRYB_31__19_), .S(SUMB_31__19_) );
  AD1V2C_8TH40 S4_20 ( .A(ab_31__20_), .B(CARRYB_30__20_), .CI(SUMB_30__21_), 
        .CO(CARRYB_31__20_), .S(SUMB_31__20_) );
  AD1V2C_8TH40 S4_21 ( .A(ab_31__21_), .B(CARRYB_30__21_), .CI(SUMB_30__22_), 
        .CO(CARRYB_31__21_), .S(SUMB_31__21_) );
  AD1V2C_8TH40 S4_22 ( .A(ab_31__22_), .B(CARRYB_30__22_), .CI(SUMB_30__23_), 
        .CO(CARRYB_31__22_), .S(SUMB_31__22_) );
  AD1V2C_8TH40 S4_23 ( .A(ab_31__23_), .B(CARRYB_30__23_), .CI(SUMB_30__24_), 
        .CO(CARRYB_31__23_), .S(SUMB_31__23_) );
  AD1V2C_8TH40 S4_24 ( .A(ab_31__24_), .B(CARRYB_30__24_), .CI(SUMB_30__25_), 
        .CO(CARRYB_31__24_), .S(SUMB_31__24_) );
  AD1V2C_8TH40 S4_25 ( .A(ab_31__25_), .B(CARRYB_30__25_), .CI(SUMB_30__26_), 
        .CO(CARRYB_31__25_), .S(SUMB_31__25_) );
  AD1V2C_8TH40 S4_26 ( .A(ab_31__26_), .B(CARRYB_30__26_), .CI(SUMB_30__27_), 
        .CO(CARRYB_31__26_), .S(SUMB_31__26_) );
  AD1V2C_8TH40 S4_27 ( .A(ab_31__27_), .B(CARRYB_30__27_), .CI(SUMB_30__28_), 
        .CO(CARRYB_31__27_), .S(SUMB_31__27_) );
  AD1V2C_8TH40 S4_28 ( .A(ab_31__28_), .B(CARRYB_30__28_), .CI(SUMB_30__29_), 
        .CO(CARRYB_31__28_), .S(SUMB_31__28_) );
  AD1V2C_8TH40 S4_29 ( .A(ab_31__29_), .B(CARRYB_30__29_), .CI(SUMB_30__30_), 
        .CO(CARRYB_31__29_), .S(SUMB_31__29_) );
  AD1V2C_8TH40 S5_30 ( .A(ab_31__30_), .B(CARRYB_30__30_), .CI(ab_30__31_), 
        .CO(CARRYB_31__30_), .S(SUMB_31__30_) );
  AD1V2C_8TH40 S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), 
        .CO(CARRYB_30__0_), .S(A1_28_) );
  AD1V2C_8TH40 S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), 
        .CO(CARRYB_30__1_), .S(SUMB_30__1_) );
  AD1V2C_8TH40 S2_30_2 ( .A(ab_30__2_), .B(CARRYB_29__2_), .CI(SUMB_29__3_), 
        .CO(CARRYB_30__2_), .S(SUMB_30__2_) );
  AD1V2C_8TH40 S2_30_3 ( .A(ab_30__3_), .B(CARRYB_29__3_), .CI(SUMB_29__4_), 
        .CO(CARRYB_30__3_), .S(SUMB_30__3_) );
  AD1V2C_8TH40 S2_30_4 ( .A(ab_30__4_), .B(CARRYB_29__4_), .CI(SUMB_29__5_), 
        .CO(CARRYB_30__4_), .S(SUMB_30__4_) );
  AD1V2C_8TH40 S2_30_5 ( .A(ab_30__5_), .B(CARRYB_29__5_), .CI(SUMB_29__6_), 
        .CO(CARRYB_30__5_), .S(SUMB_30__5_) );
  AD1V2C_8TH40 S2_30_6 ( .A(ab_30__6_), .B(CARRYB_29__6_), .CI(SUMB_29__7_), 
        .CO(CARRYB_30__6_), .S(SUMB_30__6_) );
  AD1V2C_8TH40 S2_30_7 ( .A(ab_30__7_), .B(CARRYB_29__7_), .CI(SUMB_29__8_), 
        .CO(CARRYB_30__7_), .S(SUMB_30__7_) );
  AD1V2C_8TH40 S2_30_8 ( .A(ab_30__8_), .B(CARRYB_29__8_), .CI(SUMB_29__9_), 
        .CO(CARRYB_30__8_), .S(SUMB_30__8_) );
  AD1V2C_8TH40 S2_30_9 ( .A(ab_30__9_), .B(CARRYB_29__9_), .CI(SUMB_29__10_), 
        .CO(CARRYB_30__9_), .S(SUMB_30__9_) );
  AD1V2C_8TH40 S2_30_10 ( .A(ab_30__10_), .B(CARRYB_29__10_), .CI(SUMB_29__11_), .CO(CARRYB_30__10_), .S(SUMB_30__10_) );
  AD1V2C_8TH40 S2_30_11 ( .A(ab_30__11_), .B(CARRYB_29__11_), .CI(SUMB_29__12_), .CO(CARRYB_30__11_), .S(SUMB_30__11_) );
  AD1V2C_8TH40 S2_30_12 ( .A(ab_30__12_), .B(CARRYB_29__12_), .CI(SUMB_29__13_), .CO(CARRYB_30__12_), .S(SUMB_30__12_) );
  AD1V2C_8TH40 S2_30_13 ( .A(ab_30__13_), .B(CARRYB_29__13_), .CI(SUMB_29__14_), .CO(CARRYB_30__13_), .S(SUMB_30__13_) );
  AD1V2C_8TH40 S2_30_14 ( .A(ab_30__14_), .B(CARRYB_29__14_), .CI(SUMB_29__15_), .CO(CARRYB_30__14_), .S(SUMB_30__14_) );
  AD1V2C_8TH40 S2_30_15 ( .A(ab_30__15_), .B(CARRYB_29__15_), .CI(SUMB_29__16_), .CO(CARRYB_30__15_), .S(SUMB_30__15_) );
  AD1V2C_8TH40 S2_30_16 ( .A(ab_30__16_), .B(CARRYB_29__16_), .CI(SUMB_29__17_), .CO(CARRYB_30__16_), .S(SUMB_30__16_) );
  AD1V2C_8TH40 S2_30_17 ( .A(ab_30__17_), .B(CARRYB_29__17_), .CI(SUMB_29__18_), .CO(CARRYB_30__17_), .S(SUMB_30__17_) );
  AD1V2C_8TH40 S2_30_18 ( .A(ab_30__18_), .B(CARRYB_29__18_), .CI(SUMB_29__19_), .CO(CARRYB_30__18_), .S(SUMB_30__18_) );
  AD1V2C_8TH40 S2_30_19 ( .A(ab_30__19_), .B(CARRYB_29__19_), .CI(SUMB_29__20_), .CO(CARRYB_30__19_), .S(SUMB_30__19_) );
  AD1V2C_8TH40 S2_30_20 ( .A(ab_30__20_), .B(CARRYB_29__20_), .CI(SUMB_29__21_), .CO(CARRYB_30__20_), .S(SUMB_30__20_) );
  AD1V2C_8TH40 S2_30_21 ( .A(ab_30__21_), .B(CARRYB_29__21_), .CI(SUMB_29__22_), .CO(CARRYB_30__21_), .S(SUMB_30__21_) );
  AD1V2C_8TH40 S2_30_22 ( .A(ab_30__22_), .B(CARRYB_29__22_), .CI(SUMB_29__23_), .CO(CARRYB_30__22_), .S(SUMB_30__22_) );
  AD1V2C_8TH40 S2_30_23 ( .A(ab_30__23_), .B(CARRYB_29__23_), .CI(SUMB_29__24_), .CO(CARRYB_30__23_), .S(SUMB_30__23_) );
  AD1V2C_8TH40 S2_30_24 ( .A(ab_30__24_), .B(CARRYB_29__24_), .CI(SUMB_29__25_), .CO(CARRYB_30__24_), .S(SUMB_30__24_) );
  AD1V2C_8TH40 S2_30_25 ( .A(ab_30__25_), .B(CARRYB_29__25_), .CI(SUMB_29__26_), .CO(CARRYB_30__25_), .S(SUMB_30__25_) );
  AD1V2C_8TH40 S2_30_26 ( .A(ab_30__26_), .B(CARRYB_29__26_), .CI(SUMB_29__27_), .CO(CARRYB_30__26_), .S(SUMB_30__26_) );
  AD1V2C_8TH40 S2_30_27 ( .A(ab_30__27_), .B(CARRYB_29__27_), .CI(SUMB_29__28_), .CO(CARRYB_30__27_), .S(SUMB_30__27_) );
  AD1V2C_8TH40 S2_30_28 ( .A(ab_30__28_), .B(CARRYB_29__28_), .CI(SUMB_29__29_), .CO(CARRYB_30__28_), .S(SUMB_30__28_) );
  AD1V2C_8TH40 S2_30_29 ( .A(ab_30__29_), .B(CARRYB_29__29_), .CI(SUMB_29__30_), .CO(CARRYB_30__29_), .S(SUMB_30__29_) );
  AD1V2C_8TH40 S3_30_30 ( .A(ab_30__30_), .B(CARRYB_29__30_), .CI(ab_29__31_), 
        .CO(CARRYB_30__30_), .S(SUMB_30__30_) );
  AD1V2C_8TH40 S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), 
        .CO(CARRYB_29__0_), .S(A1_27_) );
  AD1V2C_8TH40 S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), 
        .CO(CARRYB_29__1_), .S(SUMB_29__1_) );
  AD1V2C_8TH40 S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), 
        .CO(CARRYB_29__2_), .S(SUMB_29__2_) );
  AD1V2C_8TH40 S2_29_3 ( .A(ab_29__3_), .B(CARRYB_28__3_), .CI(SUMB_28__4_), 
        .CO(CARRYB_29__3_), .S(SUMB_29__3_) );
  AD1V2C_8TH40 S2_29_4 ( .A(ab_29__4_), .B(CARRYB_28__4_), .CI(SUMB_28__5_), 
        .CO(CARRYB_29__4_), .S(SUMB_29__4_) );
  AD1V2C_8TH40 S2_29_5 ( .A(ab_29__5_), .B(CARRYB_28__5_), .CI(SUMB_28__6_), 
        .CO(CARRYB_29__5_), .S(SUMB_29__5_) );
  AD1V2C_8TH40 S2_29_6 ( .A(ab_29__6_), .B(CARRYB_28__6_), .CI(SUMB_28__7_), 
        .CO(CARRYB_29__6_), .S(SUMB_29__6_) );
  AD1V2C_8TH40 S2_29_7 ( .A(ab_29__7_), .B(CARRYB_28__7_), .CI(SUMB_28__8_), 
        .CO(CARRYB_29__7_), .S(SUMB_29__7_) );
  AD1V2C_8TH40 S2_29_8 ( .A(ab_29__8_), .B(CARRYB_28__8_), .CI(SUMB_28__9_), 
        .CO(CARRYB_29__8_), .S(SUMB_29__8_) );
  AD1V2C_8TH40 S2_29_9 ( .A(ab_29__9_), .B(CARRYB_28__9_), .CI(SUMB_28__10_), 
        .CO(CARRYB_29__9_), .S(SUMB_29__9_) );
  AD1V2C_8TH40 S2_29_10 ( .A(ab_29__10_), .B(CARRYB_28__10_), .CI(SUMB_28__11_), .CO(CARRYB_29__10_), .S(SUMB_29__10_) );
  AD1V2C_8TH40 S2_29_11 ( .A(ab_29__11_), .B(CARRYB_28__11_), .CI(SUMB_28__12_), .CO(CARRYB_29__11_), .S(SUMB_29__11_) );
  AD1V2C_8TH40 S2_29_12 ( .A(ab_29__12_), .B(CARRYB_28__12_), .CI(SUMB_28__13_), .CO(CARRYB_29__12_), .S(SUMB_29__12_) );
  AD1V2C_8TH40 S2_29_13 ( .A(ab_29__13_), .B(CARRYB_28__13_), .CI(SUMB_28__14_), .CO(CARRYB_29__13_), .S(SUMB_29__13_) );
  AD1V2C_8TH40 S2_29_14 ( .A(ab_29__14_), .B(CARRYB_28__14_), .CI(SUMB_28__15_), .CO(CARRYB_29__14_), .S(SUMB_29__14_) );
  AD1V2C_8TH40 S2_29_15 ( .A(ab_29__15_), .B(CARRYB_28__15_), .CI(SUMB_28__16_), .CO(CARRYB_29__15_), .S(SUMB_29__15_) );
  AD1V2C_8TH40 S2_29_16 ( .A(ab_29__16_), .B(CARRYB_28__16_), .CI(SUMB_28__17_), .CO(CARRYB_29__16_), .S(SUMB_29__16_) );
  AD1V2C_8TH40 S2_29_17 ( .A(ab_29__17_), .B(CARRYB_28__17_), .CI(SUMB_28__18_), .CO(CARRYB_29__17_), .S(SUMB_29__17_) );
  AD1V2C_8TH40 S2_29_18 ( .A(ab_29__18_), .B(CARRYB_28__18_), .CI(SUMB_28__19_), .CO(CARRYB_29__18_), .S(SUMB_29__18_) );
  AD1V2C_8TH40 S2_29_19 ( .A(ab_29__19_), .B(CARRYB_28__19_), .CI(SUMB_28__20_), .CO(CARRYB_29__19_), .S(SUMB_29__19_) );
  AD1V2C_8TH40 S2_29_20 ( .A(ab_29__20_), .B(CARRYB_28__20_), .CI(SUMB_28__21_), .CO(CARRYB_29__20_), .S(SUMB_29__20_) );
  AD1V2C_8TH40 S2_29_21 ( .A(ab_29__21_), .B(CARRYB_28__21_), .CI(SUMB_28__22_), .CO(CARRYB_29__21_), .S(SUMB_29__21_) );
  AD1V2C_8TH40 S2_29_22 ( .A(ab_29__22_), .B(CARRYB_28__22_), .CI(SUMB_28__23_), .CO(CARRYB_29__22_), .S(SUMB_29__22_) );
  AD1V2C_8TH40 S2_29_23 ( .A(ab_29__23_), .B(CARRYB_28__23_), .CI(SUMB_28__24_), .CO(CARRYB_29__23_), .S(SUMB_29__23_) );
  AD1V2C_8TH40 S2_29_24 ( .A(ab_29__24_), .B(CARRYB_28__24_), .CI(SUMB_28__25_), .CO(CARRYB_29__24_), .S(SUMB_29__24_) );
  AD1V2C_8TH40 S2_29_25 ( .A(ab_29__25_), .B(CARRYB_28__25_), .CI(SUMB_28__26_), .CO(CARRYB_29__25_), .S(SUMB_29__25_) );
  AD1V2C_8TH40 S2_29_26 ( .A(ab_29__26_), .B(CARRYB_28__26_), .CI(SUMB_28__27_), .CO(CARRYB_29__26_), .S(SUMB_29__26_) );
  AD1V2C_8TH40 S2_29_27 ( .A(ab_29__27_), .B(CARRYB_28__27_), .CI(SUMB_28__28_), .CO(CARRYB_29__27_), .S(SUMB_29__27_) );
  AD1V2C_8TH40 S2_29_28 ( .A(ab_29__28_), .B(CARRYB_28__28_), .CI(SUMB_28__29_), .CO(CARRYB_29__28_), .S(SUMB_29__28_) );
  AD1V2C_8TH40 S2_29_29 ( .A(ab_29__29_), .B(CARRYB_28__29_), .CI(SUMB_28__30_), .CO(CARRYB_29__29_), .S(SUMB_29__29_) );
  AD1V2C_8TH40 S3_29_30 ( .A(ab_29__30_), .B(CARRYB_28__30_), .CI(ab_28__31_), 
        .CO(CARRYB_29__30_), .S(SUMB_29__30_) );
  AD1V2C_8TH40 S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), 
        .CO(CARRYB_28__0_), .S(A1_26_) );
  AD1V2C_8TH40 S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), 
        .CO(CARRYB_28__1_), .S(SUMB_28__1_) );
  AD1V2C_8TH40 S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), 
        .CO(CARRYB_28__2_), .S(SUMB_28__2_) );
  AD1V2C_8TH40 S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), 
        .CO(CARRYB_28__3_), .S(SUMB_28__3_) );
  AD1V2C_8TH40 S2_28_4 ( .A(ab_28__4_), .B(CARRYB_27__4_), .CI(SUMB_27__5_), 
        .CO(CARRYB_28__4_), .S(SUMB_28__4_) );
  AD1V2C_8TH40 S2_28_5 ( .A(ab_28__5_), .B(CARRYB_27__5_), .CI(SUMB_27__6_), 
        .CO(CARRYB_28__5_), .S(SUMB_28__5_) );
  AD1V2C_8TH40 S2_28_6 ( .A(ab_28__6_), .B(CARRYB_27__6_), .CI(SUMB_27__7_), 
        .CO(CARRYB_28__6_), .S(SUMB_28__6_) );
  AD1V2C_8TH40 S2_28_7 ( .A(ab_28__7_), .B(CARRYB_27__7_), .CI(SUMB_27__8_), 
        .CO(CARRYB_28__7_), .S(SUMB_28__7_) );
  AD1V2C_8TH40 S2_28_8 ( .A(ab_28__8_), .B(CARRYB_27__8_), .CI(SUMB_27__9_), 
        .CO(CARRYB_28__8_), .S(SUMB_28__8_) );
  AD1V2C_8TH40 S2_28_9 ( .A(ab_28__9_), .B(CARRYB_27__9_), .CI(SUMB_27__10_), 
        .CO(CARRYB_28__9_), .S(SUMB_28__9_) );
  AD1V2C_8TH40 S2_28_10 ( .A(ab_28__10_), .B(CARRYB_27__10_), .CI(SUMB_27__11_), .CO(CARRYB_28__10_), .S(SUMB_28__10_) );
  AD1V2C_8TH40 S2_28_11 ( .A(ab_28__11_), .B(CARRYB_27__11_), .CI(SUMB_27__12_), .CO(CARRYB_28__11_), .S(SUMB_28__11_) );
  AD1V2C_8TH40 S2_28_12 ( .A(ab_28__12_), .B(CARRYB_27__12_), .CI(SUMB_27__13_), .CO(CARRYB_28__12_), .S(SUMB_28__12_) );
  AD1V2C_8TH40 S2_28_13 ( .A(ab_28__13_), .B(CARRYB_27__13_), .CI(SUMB_27__14_), .CO(CARRYB_28__13_), .S(SUMB_28__13_) );
  AD1V2C_8TH40 S2_28_14 ( .A(ab_28__14_), .B(CARRYB_27__14_), .CI(SUMB_27__15_), .CO(CARRYB_28__14_), .S(SUMB_28__14_) );
  AD1V2C_8TH40 S2_28_15 ( .A(ab_28__15_), .B(CARRYB_27__15_), .CI(SUMB_27__16_), .CO(CARRYB_28__15_), .S(SUMB_28__15_) );
  AD1V2C_8TH40 S2_28_16 ( .A(ab_28__16_), .B(CARRYB_27__16_), .CI(SUMB_27__17_), .CO(CARRYB_28__16_), .S(SUMB_28__16_) );
  AD1V2C_8TH40 S2_28_17 ( .A(ab_28__17_), .B(CARRYB_27__17_), .CI(SUMB_27__18_), .CO(CARRYB_28__17_), .S(SUMB_28__17_) );
  AD1V2C_8TH40 S2_28_18 ( .A(ab_28__18_), .B(CARRYB_27__18_), .CI(SUMB_27__19_), .CO(CARRYB_28__18_), .S(SUMB_28__18_) );
  AD1V2C_8TH40 S2_28_19 ( .A(ab_28__19_), .B(CARRYB_27__19_), .CI(SUMB_27__20_), .CO(CARRYB_28__19_), .S(SUMB_28__19_) );
  AD1V2C_8TH40 S2_28_20 ( .A(ab_28__20_), .B(CARRYB_27__20_), .CI(SUMB_27__21_), .CO(CARRYB_28__20_), .S(SUMB_28__20_) );
  AD1V2C_8TH40 S2_28_21 ( .A(ab_28__21_), .B(CARRYB_27__21_), .CI(SUMB_27__22_), .CO(CARRYB_28__21_), .S(SUMB_28__21_) );
  AD1V2C_8TH40 S2_28_22 ( .A(ab_28__22_), .B(CARRYB_27__22_), .CI(SUMB_27__23_), .CO(CARRYB_28__22_), .S(SUMB_28__22_) );
  AD1V2C_8TH40 S2_28_23 ( .A(ab_28__23_), .B(CARRYB_27__23_), .CI(SUMB_27__24_), .CO(CARRYB_28__23_), .S(SUMB_28__23_) );
  AD1V2C_8TH40 S2_28_24 ( .A(ab_28__24_), .B(CARRYB_27__24_), .CI(SUMB_27__25_), .CO(CARRYB_28__24_), .S(SUMB_28__24_) );
  AD1V2C_8TH40 S2_28_25 ( .A(ab_28__25_), .B(CARRYB_27__25_), .CI(SUMB_27__26_), .CO(CARRYB_28__25_), .S(SUMB_28__25_) );
  AD1V2C_8TH40 S2_28_26 ( .A(ab_28__26_), .B(CARRYB_27__26_), .CI(SUMB_27__27_), .CO(CARRYB_28__26_), .S(SUMB_28__26_) );
  AD1V2C_8TH40 S2_28_27 ( .A(ab_28__27_), .B(CARRYB_27__27_), .CI(SUMB_27__28_), .CO(CARRYB_28__27_), .S(SUMB_28__27_) );
  AD1V2C_8TH40 S2_28_28 ( .A(ab_28__28_), .B(CARRYB_27__28_), .CI(SUMB_27__29_), .CO(CARRYB_28__28_), .S(SUMB_28__28_) );
  AD1V2C_8TH40 S2_28_29 ( .A(ab_28__29_), .B(CARRYB_27__29_), .CI(SUMB_27__30_), .CO(CARRYB_28__29_), .S(SUMB_28__29_) );
  AD1V2C_8TH40 S3_28_30 ( .A(ab_28__30_), .B(CARRYB_27__30_), .CI(ab_27__31_), 
        .CO(CARRYB_28__30_), .S(SUMB_28__30_) );
  AD1V2C_8TH40 S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), 
        .CO(CARRYB_27__0_), .S(A1_25_) );
  AD1V2C_8TH40 S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), 
        .CO(CARRYB_27__1_), .S(SUMB_27__1_) );
  AD1V2C_8TH40 S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), 
        .CO(CARRYB_27__2_), .S(SUMB_27__2_) );
  AD1V2C_8TH40 S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), 
        .CO(CARRYB_27__3_), .S(SUMB_27__3_) );
  AD1V2C_8TH40 S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), 
        .CO(CARRYB_27__4_), .S(SUMB_27__4_) );
  AD1V2C_8TH40 S2_27_5 ( .A(ab_27__5_), .B(CARRYB_26__5_), .CI(SUMB_26__6_), 
        .CO(CARRYB_27__5_), .S(SUMB_27__5_) );
  AD1V2C_8TH40 S2_27_6 ( .A(ab_27__6_), .B(CARRYB_26__6_), .CI(SUMB_26__7_), 
        .CO(CARRYB_27__6_), .S(SUMB_27__6_) );
  AD1V2C_8TH40 S2_27_7 ( .A(ab_27__7_), .B(CARRYB_26__7_), .CI(SUMB_26__8_), 
        .CO(CARRYB_27__7_), .S(SUMB_27__7_) );
  AD1V2C_8TH40 S2_27_8 ( .A(ab_27__8_), .B(CARRYB_26__8_), .CI(SUMB_26__9_), 
        .CO(CARRYB_27__8_), .S(SUMB_27__8_) );
  AD1V2C_8TH40 S2_27_9 ( .A(ab_27__9_), .B(CARRYB_26__9_), .CI(SUMB_26__10_), 
        .CO(CARRYB_27__9_), .S(SUMB_27__9_) );
  AD1V2C_8TH40 S2_27_10 ( .A(ab_27__10_), .B(CARRYB_26__10_), .CI(SUMB_26__11_), .CO(CARRYB_27__10_), .S(SUMB_27__10_) );
  AD1V2C_8TH40 S2_27_11 ( .A(ab_27__11_), .B(CARRYB_26__11_), .CI(SUMB_26__12_), .CO(CARRYB_27__11_), .S(SUMB_27__11_) );
  AD1V2C_8TH40 S2_27_12 ( .A(ab_27__12_), .B(CARRYB_26__12_), .CI(SUMB_26__13_), .CO(CARRYB_27__12_), .S(SUMB_27__12_) );
  AD1V2C_8TH40 S2_27_13 ( .A(ab_27__13_), .B(CARRYB_26__13_), .CI(SUMB_26__14_), .CO(CARRYB_27__13_), .S(SUMB_27__13_) );
  AD1V2C_8TH40 S2_27_14 ( .A(ab_27__14_), .B(CARRYB_26__14_), .CI(SUMB_26__15_), .CO(CARRYB_27__14_), .S(SUMB_27__14_) );
  AD1V2C_8TH40 S2_27_15 ( .A(ab_27__15_), .B(CARRYB_26__15_), .CI(SUMB_26__16_), .CO(CARRYB_27__15_), .S(SUMB_27__15_) );
  AD1V2C_8TH40 S2_27_16 ( .A(ab_27__16_), .B(CARRYB_26__16_), .CI(SUMB_26__17_), .CO(CARRYB_27__16_), .S(SUMB_27__16_) );
  AD1V2C_8TH40 S2_27_17 ( .A(ab_27__17_), .B(CARRYB_26__17_), .CI(SUMB_26__18_), .CO(CARRYB_27__17_), .S(SUMB_27__17_) );
  AD1V2C_8TH40 S2_27_18 ( .A(ab_27__18_), .B(CARRYB_26__18_), .CI(SUMB_26__19_), .CO(CARRYB_27__18_), .S(SUMB_27__18_) );
  AD1V2C_8TH40 S2_27_19 ( .A(ab_27__19_), .B(CARRYB_26__19_), .CI(SUMB_26__20_), .CO(CARRYB_27__19_), .S(SUMB_27__19_) );
  AD1V2C_8TH40 S2_27_20 ( .A(ab_27__20_), .B(CARRYB_26__20_), .CI(SUMB_26__21_), .CO(CARRYB_27__20_), .S(SUMB_27__20_) );
  AD1V2C_8TH40 S2_27_21 ( .A(ab_27__21_), .B(CARRYB_26__21_), .CI(SUMB_26__22_), .CO(CARRYB_27__21_), .S(SUMB_27__21_) );
  AD1V2C_8TH40 S2_27_22 ( .A(ab_27__22_), .B(CARRYB_26__22_), .CI(SUMB_26__23_), .CO(CARRYB_27__22_), .S(SUMB_27__22_) );
  AD1V2C_8TH40 S2_27_23 ( .A(ab_27__23_), .B(CARRYB_26__23_), .CI(SUMB_26__24_), .CO(CARRYB_27__23_), .S(SUMB_27__23_) );
  AD1V2C_8TH40 S2_27_24 ( .A(ab_27__24_), .B(CARRYB_26__24_), .CI(SUMB_26__25_), .CO(CARRYB_27__24_), .S(SUMB_27__24_) );
  AD1V2C_8TH40 S2_27_25 ( .A(ab_27__25_), .B(CARRYB_26__25_), .CI(SUMB_26__26_), .CO(CARRYB_27__25_), .S(SUMB_27__25_) );
  AD1V2C_8TH40 S2_27_26 ( .A(ab_27__26_), .B(CARRYB_26__26_), .CI(SUMB_26__27_), .CO(CARRYB_27__26_), .S(SUMB_27__26_) );
  AD1V2C_8TH40 S2_27_27 ( .A(ab_27__27_), .B(CARRYB_26__27_), .CI(SUMB_26__28_), .CO(CARRYB_27__27_), .S(SUMB_27__27_) );
  AD1V2C_8TH40 S2_27_28 ( .A(ab_27__28_), .B(CARRYB_26__28_), .CI(SUMB_26__29_), .CO(CARRYB_27__28_), .S(SUMB_27__28_) );
  AD1V2C_8TH40 S2_27_29 ( .A(ab_27__29_), .B(CARRYB_26__29_), .CI(SUMB_26__30_), .CO(CARRYB_27__29_), .S(SUMB_27__29_) );
  AD1V2C_8TH40 S3_27_30 ( .A(ab_27__30_), .B(CARRYB_26__30_), .CI(ab_26__31_), 
        .CO(CARRYB_27__30_), .S(SUMB_27__30_) );
  AD1V2C_8TH40 S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), 
        .CO(CARRYB_26__0_), .S(A1_24_) );
  AD1V2C_8TH40 S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), 
        .CO(CARRYB_26__1_), .S(SUMB_26__1_) );
  AD1V2C_8TH40 S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), 
        .CO(CARRYB_26__2_), .S(SUMB_26__2_) );
  AD1V2C_8TH40 S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), 
        .CO(CARRYB_26__3_), .S(SUMB_26__3_) );
  AD1V2C_8TH40 S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), 
        .CO(CARRYB_26__4_), .S(SUMB_26__4_) );
  AD1V2C_8TH40 S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), 
        .CO(CARRYB_26__5_), .S(SUMB_26__5_) );
  AD1V2C_8TH40 S2_26_6 ( .A(ab_26__6_), .B(CARRYB_25__6_), .CI(SUMB_25__7_), 
        .CO(CARRYB_26__6_), .S(SUMB_26__6_) );
  AD1V2C_8TH40 S2_26_7 ( .A(ab_26__7_), .B(CARRYB_25__7_), .CI(SUMB_25__8_), 
        .CO(CARRYB_26__7_), .S(SUMB_26__7_) );
  AD1V2C_8TH40 S2_26_8 ( .A(ab_26__8_), .B(CARRYB_25__8_), .CI(SUMB_25__9_), 
        .CO(CARRYB_26__8_), .S(SUMB_26__8_) );
  AD1V2C_8TH40 S2_26_9 ( .A(ab_26__9_), .B(CARRYB_25__9_), .CI(SUMB_25__10_), 
        .CO(CARRYB_26__9_), .S(SUMB_26__9_) );
  AD1V2C_8TH40 S2_26_10 ( .A(ab_26__10_), .B(CARRYB_25__10_), .CI(SUMB_25__11_), .CO(CARRYB_26__10_), .S(SUMB_26__10_) );
  AD1V2C_8TH40 S2_26_11 ( .A(ab_26__11_), .B(CARRYB_25__11_), .CI(SUMB_25__12_), .CO(CARRYB_26__11_), .S(SUMB_26__11_) );
  AD1V2C_8TH40 S2_26_12 ( .A(ab_26__12_), .B(CARRYB_25__12_), .CI(SUMB_25__13_), .CO(CARRYB_26__12_), .S(SUMB_26__12_) );
  AD1V2C_8TH40 S2_26_13 ( .A(ab_26__13_), .B(CARRYB_25__13_), .CI(SUMB_25__14_), .CO(CARRYB_26__13_), .S(SUMB_26__13_) );
  AD1V2C_8TH40 S2_26_14 ( .A(ab_26__14_), .B(CARRYB_25__14_), .CI(SUMB_25__15_), .CO(CARRYB_26__14_), .S(SUMB_26__14_) );
  AD1V2C_8TH40 S2_26_15 ( .A(ab_26__15_), .B(CARRYB_25__15_), .CI(SUMB_25__16_), .CO(CARRYB_26__15_), .S(SUMB_26__15_) );
  AD1V2C_8TH40 S2_26_16 ( .A(ab_26__16_), .B(CARRYB_25__16_), .CI(SUMB_25__17_), .CO(CARRYB_26__16_), .S(SUMB_26__16_) );
  AD1V2C_8TH40 S2_26_17 ( .A(ab_26__17_), .B(CARRYB_25__17_), .CI(SUMB_25__18_), .CO(CARRYB_26__17_), .S(SUMB_26__17_) );
  AD1V2C_8TH40 S2_26_18 ( .A(ab_26__18_), .B(CARRYB_25__18_), .CI(SUMB_25__19_), .CO(CARRYB_26__18_), .S(SUMB_26__18_) );
  AD1V2C_8TH40 S2_26_19 ( .A(ab_26__19_), .B(CARRYB_25__19_), .CI(SUMB_25__20_), .CO(CARRYB_26__19_), .S(SUMB_26__19_) );
  AD1V2C_8TH40 S2_26_20 ( .A(ab_26__20_), .B(CARRYB_25__20_), .CI(SUMB_25__21_), .CO(CARRYB_26__20_), .S(SUMB_26__20_) );
  AD1V2C_8TH40 S2_26_21 ( .A(ab_26__21_), .B(CARRYB_25__21_), .CI(SUMB_25__22_), .CO(CARRYB_26__21_), .S(SUMB_26__21_) );
  AD1V2C_8TH40 S2_26_22 ( .A(ab_26__22_), .B(CARRYB_25__22_), .CI(SUMB_25__23_), .CO(CARRYB_26__22_), .S(SUMB_26__22_) );
  AD1V2C_8TH40 S2_26_23 ( .A(ab_26__23_), .B(CARRYB_25__23_), .CI(SUMB_25__24_), .CO(CARRYB_26__23_), .S(SUMB_26__23_) );
  AD1V2C_8TH40 S2_26_24 ( .A(ab_26__24_), .B(CARRYB_25__24_), .CI(SUMB_25__25_), .CO(CARRYB_26__24_), .S(SUMB_26__24_) );
  AD1V2C_8TH40 S2_26_25 ( .A(ab_26__25_), .B(CARRYB_25__25_), .CI(SUMB_25__26_), .CO(CARRYB_26__25_), .S(SUMB_26__25_) );
  AD1V2C_8TH40 S2_26_26 ( .A(ab_26__26_), .B(CARRYB_25__26_), .CI(SUMB_25__27_), .CO(CARRYB_26__26_), .S(SUMB_26__26_) );
  AD1V2C_8TH40 S2_26_27 ( .A(ab_26__27_), .B(CARRYB_25__27_), .CI(SUMB_25__28_), .CO(CARRYB_26__27_), .S(SUMB_26__27_) );
  AD1V2C_8TH40 S2_26_28 ( .A(ab_26__28_), .B(CARRYB_25__28_), .CI(SUMB_25__29_), .CO(CARRYB_26__28_), .S(SUMB_26__28_) );
  AD1V2C_8TH40 S2_26_29 ( .A(ab_26__29_), .B(CARRYB_25__29_), .CI(SUMB_25__30_), .CO(CARRYB_26__29_), .S(SUMB_26__29_) );
  AD1V2C_8TH40 S3_26_30 ( .A(ab_26__30_), .B(CARRYB_25__30_), .CI(ab_25__31_), 
        .CO(CARRYB_26__30_), .S(SUMB_26__30_) );
  AD1V2C_8TH40 S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), 
        .CO(CARRYB_25__0_), .S(A1_23_) );
  AD1V2C_8TH40 S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), 
        .CO(CARRYB_25__1_), .S(SUMB_25__1_) );
  AD1V2C_8TH40 S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), 
        .CO(CARRYB_25__2_), .S(SUMB_25__2_) );
  AD1V2C_8TH40 S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), 
        .CO(CARRYB_25__3_), .S(SUMB_25__3_) );
  AD1V2C_8TH40 S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), 
        .CO(CARRYB_25__4_), .S(SUMB_25__4_) );
  AD1V2C_8TH40 S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), 
        .CO(CARRYB_25__5_), .S(SUMB_25__5_) );
  AD1V2C_8TH40 S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), 
        .CO(CARRYB_25__6_), .S(SUMB_25__6_) );
  AD1V2C_8TH40 S2_25_7 ( .A(ab_25__7_), .B(CARRYB_24__7_), .CI(SUMB_24__8_), 
        .CO(CARRYB_25__7_), .S(SUMB_25__7_) );
  AD1V2C_8TH40 S2_25_8 ( .A(ab_25__8_), .B(CARRYB_24__8_), .CI(SUMB_24__9_), 
        .CO(CARRYB_25__8_), .S(SUMB_25__8_) );
  AD1V2C_8TH40 S2_25_9 ( .A(ab_25__9_), .B(CARRYB_24__9_), .CI(SUMB_24__10_), 
        .CO(CARRYB_25__9_), .S(SUMB_25__9_) );
  AD1V2C_8TH40 S2_25_10 ( .A(ab_25__10_), .B(CARRYB_24__10_), .CI(SUMB_24__11_), .CO(CARRYB_25__10_), .S(SUMB_25__10_) );
  AD1V2C_8TH40 S2_25_11 ( .A(ab_25__11_), .B(CARRYB_24__11_), .CI(SUMB_24__12_), .CO(CARRYB_25__11_), .S(SUMB_25__11_) );
  AD1V2C_8TH40 S2_25_12 ( .A(ab_25__12_), .B(CARRYB_24__12_), .CI(SUMB_24__13_), .CO(CARRYB_25__12_), .S(SUMB_25__12_) );
  AD1V2C_8TH40 S2_25_13 ( .A(ab_25__13_), .B(CARRYB_24__13_), .CI(SUMB_24__14_), .CO(CARRYB_25__13_), .S(SUMB_25__13_) );
  AD1V2C_8TH40 S2_25_14 ( .A(ab_25__14_), .B(CARRYB_24__14_), .CI(SUMB_24__15_), .CO(CARRYB_25__14_), .S(SUMB_25__14_) );
  AD1V2C_8TH40 S2_25_15 ( .A(ab_25__15_), .B(CARRYB_24__15_), .CI(SUMB_24__16_), .CO(CARRYB_25__15_), .S(SUMB_25__15_) );
  AD1V2C_8TH40 S2_25_16 ( .A(ab_25__16_), .B(CARRYB_24__16_), .CI(SUMB_24__17_), .CO(CARRYB_25__16_), .S(SUMB_25__16_) );
  AD1V2C_8TH40 S2_25_17 ( .A(ab_25__17_), .B(CARRYB_24__17_), .CI(SUMB_24__18_), .CO(CARRYB_25__17_), .S(SUMB_25__17_) );
  AD1V2C_8TH40 S2_25_18 ( .A(ab_25__18_), .B(CARRYB_24__18_), .CI(SUMB_24__19_), .CO(CARRYB_25__18_), .S(SUMB_25__18_) );
  AD1V2C_8TH40 S2_25_19 ( .A(ab_25__19_), .B(CARRYB_24__19_), .CI(SUMB_24__20_), .CO(CARRYB_25__19_), .S(SUMB_25__19_) );
  AD1V2C_8TH40 S2_25_20 ( .A(ab_25__20_), .B(CARRYB_24__20_), .CI(SUMB_24__21_), .CO(CARRYB_25__20_), .S(SUMB_25__20_) );
  AD1V2C_8TH40 S2_25_21 ( .A(ab_25__21_), .B(CARRYB_24__21_), .CI(SUMB_24__22_), .CO(CARRYB_25__21_), .S(SUMB_25__21_) );
  AD1V2C_8TH40 S2_25_22 ( .A(ab_25__22_), .B(CARRYB_24__22_), .CI(SUMB_24__23_), .CO(CARRYB_25__22_), .S(SUMB_25__22_) );
  AD1V2C_8TH40 S2_25_23 ( .A(ab_25__23_), .B(CARRYB_24__23_), .CI(SUMB_24__24_), .CO(CARRYB_25__23_), .S(SUMB_25__23_) );
  AD1V2C_8TH40 S2_25_24 ( .A(ab_25__24_), .B(CARRYB_24__24_), .CI(SUMB_24__25_), .CO(CARRYB_25__24_), .S(SUMB_25__24_) );
  AD1V2C_8TH40 S2_25_25 ( .A(ab_25__25_), .B(CARRYB_24__25_), .CI(SUMB_24__26_), .CO(CARRYB_25__25_), .S(SUMB_25__25_) );
  AD1V2C_8TH40 S2_25_26 ( .A(ab_25__26_), .B(CARRYB_24__26_), .CI(SUMB_24__27_), .CO(CARRYB_25__26_), .S(SUMB_25__26_) );
  AD1V2C_8TH40 S2_25_27 ( .A(ab_25__27_), .B(CARRYB_24__27_), .CI(SUMB_24__28_), .CO(CARRYB_25__27_), .S(SUMB_25__27_) );
  AD1V2C_8TH40 S2_25_28 ( .A(ab_25__28_), .B(CARRYB_24__28_), .CI(SUMB_24__29_), .CO(CARRYB_25__28_), .S(SUMB_25__28_) );
  AD1V2C_8TH40 S2_25_29 ( .A(ab_25__29_), .B(CARRYB_24__29_), .CI(SUMB_24__30_), .CO(CARRYB_25__29_), .S(SUMB_25__29_) );
  AD1V2C_8TH40 S3_25_30 ( .A(ab_25__30_), .B(CARRYB_24__30_), .CI(ab_24__31_), 
        .CO(CARRYB_25__30_), .S(SUMB_25__30_) );
  AD1V2C_8TH40 S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), 
        .CO(CARRYB_24__0_), .S(A1_22_) );
  AD1V2C_8TH40 S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), 
        .CO(CARRYB_24__1_), .S(SUMB_24__1_) );
  AD1V2C_8TH40 S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), 
        .CO(CARRYB_24__2_), .S(SUMB_24__2_) );
  AD1V2C_8TH40 S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), 
        .CO(CARRYB_24__3_), .S(SUMB_24__3_) );
  AD1V2C_8TH40 S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), 
        .CO(CARRYB_24__4_), .S(SUMB_24__4_) );
  AD1V2C_8TH40 S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), 
        .CO(CARRYB_24__5_), .S(SUMB_24__5_) );
  AD1V2C_8TH40 S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), 
        .CO(CARRYB_24__6_), .S(SUMB_24__6_) );
  AD1V2C_8TH40 S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), 
        .CO(CARRYB_24__7_), .S(SUMB_24__7_) );
  AD1V2C_8TH40 S2_24_8 ( .A(ab_24__8_), .B(CARRYB_23__8_), .CI(SUMB_23__9_), 
        .CO(CARRYB_24__8_), .S(SUMB_24__8_) );
  AD1V2C_8TH40 S2_24_9 ( .A(ab_24__9_), .B(CARRYB_23__9_), .CI(SUMB_23__10_), 
        .CO(CARRYB_24__9_), .S(SUMB_24__9_) );
  AD1V2C_8TH40 S2_24_10 ( .A(ab_24__10_), .B(CARRYB_23__10_), .CI(SUMB_23__11_), .CO(CARRYB_24__10_), .S(SUMB_24__10_) );
  AD1V2C_8TH40 S2_24_11 ( .A(ab_24__11_), .B(CARRYB_23__11_), .CI(SUMB_23__12_), .CO(CARRYB_24__11_), .S(SUMB_24__11_) );
  AD1V2C_8TH40 S2_24_12 ( .A(ab_24__12_), .B(CARRYB_23__12_), .CI(SUMB_23__13_), .CO(CARRYB_24__12_), .S(SUMB_24__12_) );
  AD1V2C_8TH40 S2_24_13 ( .A(ab_24__13_), .B(CARRYB_23__13_), .CI(SUMB_23__14_), .CO(CARRYB_24__13_), .S(SUMB_24__13_) );
  AD1V2C_8TH40 S2_24_14 ( .A(ab_24__14_), .B(CARRYB_23__14_), .CI(SUMB_23__15_), .CO(CARRYB_24__14_), .S(SUMB_24__14_) );
  AD1V2C_8TH40 S2_24_15 ( .A(ab_24__15_), .B(CARRYB_23__15_), .CI(SUMB_23__16_), .CO(CARRYB_24__15_), .S(SUMB_24__15_) );
  AD1V2C_8TH40 S2_24_16 ( .A(ab_24__16_), .B(CARRYB_23__16_), .CI(SUMB_23__17_), .CO(CARRYB_24__16_), .S(SUMB_24__16_) );
  AD1V2C_8TH40 S2_24_17 ( .A(ab_24__17_), .B(CARRYB_23__17_), .CI(SUMB_23__18_), .CO(CARRYB_24__17_), .S(SUMB_24__17_) );
  AD1V2C_8TH40 S2_24_18 ( .A(ab_24__18_), .B(CARRYB_23__18_), .CI(SUMB_23__19_), .CO(CARRYB_24__18_), .S(SUMB_24__18_) );
  AD1V2C_8TH40 S2_24_19 ( .A(ab_24__19_), .B(CARRYB_23__19_), .CI(SUMB_23__20_), .CO(CARRYB_24__19_), .S(SUMB_24__19_) );
  AD1V2C_8TH40 S2_24_20 ( .A(ab_24__20_), .B(CARRYB_23__20_), .CI(SUMB_23__21_), .CO(CARRYB_24__20_), .S(SUMB_24__20_) );
  AD1V2C_8TH40 S2_24_21 ( .A(ab_24__21_), .B(CARRYB_23__21_), .CI(SUMB_23__22_), .CO(CARRYB_24__21_), .S(SUMB_24__21_) );
  AD1V2C_8TH40 S2_24_22 ( .A(ab_24__22_), .B(CARRYB_23__22_), .CI(SUMB_23__23_), .CO(CARRYB_24__22_), .S(SUMB_24__22_) );
  AD1V2C_8TH40 S2_24_23 ( .A(ab_24__23_), .B(CARRYB_23__23_), .CI(SUMB_23__24_), .CO(CARRYB_24__23_), .S(SUMB_24__23_) );
  AD1V2C_8TH40 S2_24_24 ( .A(ab_24__24_), .B(CARRYB_23__24_), .CI(SUMB_23__25_), .CO(CARRYB_24__24_), .S(SUMB_24__24_) );
  AD1V2C_8TH40 S2_24_25 ( .A(ab_24__25_), .B(CARRYB_23__25_), .CI(SUMB_23__26_), .CO(CARRYB_24__25_), .S(SUMB_24__25_) );
  AD1V2C_8TH40 S2_24_26 ( .A(ab_24__26_), .B(CARRYB_23__26_), .CI(SUMB_23__27_), .CO(CARRYB_24__26_), .S(SUMB_24__26_) );
  AD1V2C_8TH40 S2_24_27 ( .A(ab_24__27_), .B(CARRYB_23__27_), .CI(SUMB_23__28_), .CO(CARRYB_24__27_), .S(SUMB_24__27_) );
  AD1V2C_8TH40 S2_24_28 ( .A(ab_24__28_), .B(CARRYB_23__28_), .CI(SUMB_23__29_), .CO(CARRYB_24__28_), .S(SUMB_24__28_) );
  AD1V2C_8TH40 S2_24_29 ( .A(ab_24__29_), .B(CARRYB_23__29_), .CI(SUMB_23__30_), .CO(CARRYB_24__29_), .S(SUMB_24__29_) );
  AD1V2C_8TH40 S3_24_30 ( .A(ab_24__30_), .B(CARRYB_23__30_), .CI(ab_23__31_), 
        .CO(CARRYB_24__30_), .S(SUMB_24__30_) );
  AD1V2C_8TH40 S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), 
        .CO(CARRYB_23__0_), .S(A1_21_) );
  AD1V2C_8TH40 S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), 
        .CO(CARRYB_23__1_), .S(SUMB_23__1_) );
  AD1V2C_8TH40 S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), 
        .CO(CARRYB_23__2_), .S(SUMB_23__2_) );
  AD1V2C_8TH40 S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), 
        .CO(CARRYB_23__3_), .S(SUMB_23__3_) );
  AD1V2C_8TH40 S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), 
        .CO(CARRYB_23__4_), .S(SUMB_23__4_) );
  AD1V2C_8TH40 S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), 
        .CO(CARRYB_23__5_), .S(SUMB_23__5_) );
  AD1V2C_8TH40 S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), 
        .CO(CARRYB_23__6_), .S(SUMB_23__6_) );
  AD1V2C_8TH40 S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), 
        .CO(CARRYB_23__7_), .S(SUMB_23__7_) );
  AD1V2C_8TH40 S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), 
        .CO(CARRYB_23__8_), .S(SUMB_23__8_) );
  AD1V2C_8TH40 S2_23_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), 
        .CO(CARRYB_23__9_), .S(SUMB_23__9_) );
  AD1V2C_8TH40 S2_23_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(CARRYB_23__10_), .S(SUMB_23__10_) );
  AD1V2C_8TH40 S2_23_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(CARRYB_23__11_), .S(SUMB_23__11_) );
  AD1V2C_8TH40 S2_23_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(CARRYB_23__12_), .S(SUMB_23__12_) );
  AD1V2C_8TH40 S2_23_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(CARRYB_23__13_), .S(SUMB_23__13_) );
  AD1V2C_8TH40 S2_23_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(CARRYB_23__14_), .S(SUMB_23__14_) );
  AD1V2C_8TH40 S2_23_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(CARRYB_23__15_), .S(SUMB_23__15_) );
  AD1V2C_8TH40 S2_23_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(CARRYB_23__16_), .S(SUMB_23__16_) );
  AD1V2C_8TH40 S2_23_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(CARRYB_23__17_), .S(SUMB_23__17_) );
  AD1V2C_8TH40 S2_23_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(CARRYB_23__18_), .S(SUMB_23__18_) );
  AD1V2C_8TH40 S2_23_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(CARRYB_23__19_), .S(SUMB_23__19_) );
  AD1V2C_8TH40 S2_23_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(CARRYB_23__20_), .S(SUMB_23__20_) );
  AD1V2C_8TH40 S2_23_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(CARRYB_23__21_), .S(SUMB_23__21_) );
  AD1V2C_8TH40 S2_23_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(SUMB_22__23_), .CO(CARRYB_23__22_), .S(SUMB_23__22_) );
  AD1V2C_8TH40 S2_23_23 ( .A(ab_23__23_), .B(CARRYB_22__23_), .CI(SUMB_22__24_), .CO(CARRYB_23__23_), .S(SUMB_23__23_) );
  AD1V2C_8TH40 S2_23_24 ( .A(ab_23__24_), .B(CARRYB_22__24_), .CI(SUMB_22__25_), .CO(CARRYB_23__24_), .S(SUMB_23__24_) );
  AD1V2C_8TH40 S2_23_25 ( .A(ab_23__25_), .B(CARRYB_22__25_), .CI(SUMB_22__26_), .CO(CARRYB_23__25_), .S(SUMB_23__25_) );
  AD1V2C_8TH40 S2_23_26 ( .A(ab_23__26_), .B(CARRYB_22__26_), .CI(SUMB_22__27_), .CO(CARRYB_23__26_), .S(SUMB_23__26_) );
  AD1V2C_8TH40 S2_23_27 ( .A(ab_23__27_), .B(CARRYB_22__27_), .CI(SUMB_22__28_), .CO(CARRYB_23__27_), .S(SUMB_23__27_) );
  AD1V2C_8TH40 S2_23_28 ( .A(ab_23__28_), .B(CARRYB_22__28_), .CI(SUMB_22__29_), .CO(CARRYB_23__28_), .S(SUMB_23__28_) );
  AD1V2C_8TH40 S2_23_29 ( .A(ab_23__29_), .B(CARRYB_22__29_), .CI(SUMB_22__30_), .CO(CARRYB_23__29_), .S(SUMB_23__29_) );
  AD1V2C_8TH40 S3_23_30 ( .A(ab_23__30_), .B(CARRYB_22__30_), .CI(ab_22__31_), 
        .CO(CARRYB_23__30_), .S(SUMB_23__30_) );
  AD1V2C_8TH40 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), 
        .CO(CARRYB_22__0_), .S(A1_20_) );
  AD1V2C_8TH40 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), 
        .CO(CARRYB_22__1_), .S(SUMB_22__1_) );
  AD1V2C_8TH40 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), 
        .CO(CARRYB_22__2_), .S(SUMB_22__2_) );
  AD1V2C_8TH40 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), 
        .CO(CARRYB_22__3_), .S(SUMB_22__3_) );
  AD1V2C_8TH40 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), 
        .CO(CARRYB_22__4_), .S(SUMB_22__4_) );
  AD1V2C_8TH40 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), 
        .CO(CARRYB_22__5_), .S(SUMB_22__5_) );
  AD1V2C_8TH40 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), 
        .CO(CARRYB_22__6_), .S(SUMB_22__6_) );
  AD1V2C_8TH40 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), 
        .CO(CARRYB_22__7_), .S(SUMB_22__7_) );
  AD1V2C_8TH40 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), 
        .CO(CARRYB_22__8_), .S(SUMB_22__8_) );
  AD1V2C_8TH40 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), 
        .CO(CARRYB_22__9_), .S(SUMB_22__9_) );
  AD1V2C_8TH40 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(CARRYB_22__10_), .S(SUMB_22__10_) );
  AD1V2C_8TH40 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(CARRYB_22__11_), .S(SUMB_22__11_) );
  AD1V2C_8TH40 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(CARRYB_22__12_), .S(SUMB_22__12_) );
  AD1V2C_8TH40 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(CARRYB_22__13_), .S(SUMB_22__13_) );
  AD1V2C_8TH40 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(CARRYB_22__14_), .S(SUMB_22__14_) );
  AD1V2C_8TH40 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(CARRYB_22__15_), .S(SUMB_22__15_) );
  AD1V2C_8TH40 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(CARRYB_22__16_), .S(SUMB_22__16_) );
  AD1V2C_8TH40 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(CARRYB_22__17_), .S(SUMB_22__17_) );
  AD1V2C_8TH40 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(CARRYB_22__18_), .S(SUMB_22__18_) );
  AD1V2C_8TH40 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(CARRYB_22__19_), .S(SUMB_22__19_) );
  AD1V2C_8TH40 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(CARRYB_22__20_), .S(SUMB_22__20_) );
  AD1V2C_8TH40 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(CARRYB_22__21_), .S(SUMB_22__21_) );
  AD1V2C_8TH40 S2_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(SUMB_21__23_), .CO(CARRYB_22__22_), .S(SUMB_22__22_) );
  AD1V2C_8TH40 S2_22_23 ( .A(ab_22__23_), .B(CARRYB_21__23_), .CI(SUMB_21__24_), .CO(CARRYB_22__23_), .S(SUMB_22__23_) );
  AD1V2C_8TH40 S2_22_24 ( .A(ab_22__24_), .B(CARRYB_21__24_), .CI(SUMB_21__25_), .CO(CARRYB_22__24_), .S(SUMB_22__24_) );
  AD1V2C_8TH40 S2_22_25 ( .A(ab_22__25_), .B(CARRYB_21__25_), .CI(SUMB_21__26_), .CO(CARRYB_22__25_), .S(SUMB_22__25_) );
  AD1V2C_8TH40 S2_22_26 ( .A(ab_22__26_), .B(CARRYB_21__26_), .CI(SUMB_21__27_), .CO(CARRYB_22__26_), .S(SUMB_22__26_) );
  AD1V2C_8TH40 S2_22_27 ( .A(ab_22__27_), .B(CARRYB_21__27_), .CI(SUMB_21__28_), .CO(CARRYB_22__27_), .S(SUMB_22__27_) );
  AD1V2C_8TH40 S2_22_28 ( .A(ab_22__28_), .B(CARRYB_21__28_), .CI(SUMB_21__29_), .CO(CARRYB_22__28_), .S(SUMB_22__28_) );
  AD1V2C_8TH40 S2_22_29 ( .A(ab_22__29_), .B(CARRYB_21__29_), .CI(SUMB_21__30_), .CO(CARRYB_22__29_), .S(SUMB_22__29_) );
  AD1V2C_8TH40 S3_22_30 ( .A(ab_22__30_), .B(CARRYB_21__30_), .CI(ab_21__31_), 
        .CO(CARRYB_22__30_), .S(SUMB_22__30_) );
  AD1V2C_8TH40 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), 
        .CO(CARRYB_21__0_), .S(A1_19_) );
  AD1V2C_8TH40 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), 
        .CO(CARRYB_21__1_), .S(SUMB_21__1_) );
  AD1V2C_8TH40 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), 
        .CO(CARRYB_21__2_), .S(SUMB_21__2_) );
  AD1V2C_8TH40 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), 
        .CO(CARRYB_21__3_), .S(SUMB_21__3_) );
  AD1V2C_8TH40 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), 
        .CO(CARRYB_21__4_), .S(SUMB_21__4_) );
  AD1V2C_8TH40 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), 
        .CO(CARRYB_21__5_), .S(SUMB_21__5_) );
  AD1V2C_8TH40 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), 
        .CO(CARRYB_21__6_), .S(SUMB_21__6_) );
  AD1V2C_8TH40 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), 
        .CO(CARRYB_21__7_), .S(SUMB_21__7_) );
  AD1V2C_8TH40 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), 
        .CO(CARRYB_21__8_), .S(SUMB_21__8_) );
  AD1V2C_8TH40 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), 
        .CO(CARRYB_21__9_), .S(SUMB_21__9_) );
  AD1V2C_8TH40 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(CARRYB_21__10_), .S(SUMB_21__10_) );
  AD1V2C_8TH40 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(CARRYB_21__11_), .S(SUMB_21__11_) );
  AD1V2C_8TH40 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(CARRYB_21__12_), .S(SUMB_21__12_) );
  AD1V2C_8TH40 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(CARRYB_21__13_), .S(SUMB_21__13_) );
  AD1V2C_8TH40 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(CARRYB_21__14_), .S(SUMB_21__14_) );
  AD1V2C_8TH40 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(CARRYB_21__15_), .S(SUMB_21__15_) );
  AD1V2C_8TH40 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(CARRYB_21__16_), .S(SUMB_21__16_) );
  AD1V2C_8TH40 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(CARRYB_21__17_), .S(SUMB_21__17_) );
  AD1V2C_8TH40 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(CARRYB_21__18_), .S(SUMB_21__18_) );
  AD1V2C_8TH40 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(CARRYB_21__19_), .S(SUMB_21__19_) );
  AD1V2C_8TH40 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(CARRYB_21__20_), .S(SUMB_21__20_) );
  AD1V2C_8TH40 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(CARRYB_21__21_), .S(SUMB_21__21_) );
  AD1V2C_8TH40 S2_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(SUMB_20__23_), .CO(CARRYB_21__22_), .S(SUMB_21__22_) );
  AD1V2C_8TH40 S2_21_23 ( .A(ab_21__23_), .B(CARRYB_20__23_), .CI(SUMB_20__24_), .CO(CARRYB_21__23_), .S(SUMB_21__23_) );
  AD1V2C_8TH40 S2_21_24 ( .A(ab_21__24_), .B(CARRYB_20__24_), .CI(SUMB_20__25_), .CO(CARRYB_21__24_), .S(SUMB_21__24_) );
  AD1V2C_8TH40 S2_21_25 ( .A(ab_21__25_), .B(CARRYB_20__25_), .CI(SUMB_20__26_), .CO(CARRYB_21__25_), .S(SUMB_21__25_) );
  AD1V2C_8TH40 S2_21_26 ( .A(ab_21__26_), .B(CARRYB_20__26_), .CI(SUMB_20__27_), .CO(CARRYB_21__26_), .S(SUMB_21__26_) );
  AD1V2C_8TH40 S2_21_27 ( .A(ab_21__27_), .B(CARRYB_20__27_), .CI(SUMB_20__28_), .CO(CARRYB_21__27_), .S(SUMB_21__27_) );
  AD1V2C_8TH40 S2_21_28 ( .A(ab_21__28_), .B(CARRYB_20__28_), .CI(SUMB_20__29_), .CO(CARRYB_21__28_), .S(SUMB_21__28_) );
  AD1V2C_8TH40 S2_21_29 ( .A(ab_21__29_), .B(CARRYB_20__29_), .CI(SUMB_20__30_), .CO(CARRYB_21__29_), .S(SUMB_21__29_) );
  AD1V2C_8TH40 S3_21_30 ( .A(ab_21__30_), .B(CARRYB_20__30_), .CI(ab_20__31_), 
        .CO(CARRYB_21__30_), .S(SUMB_21__30_) );
  AD1V2C_8TH40 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), 
        .CO(CARRYB_20__0_), .S(A1_18_) );
  AD1V2C_8TH40 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), 
        .CO(CARRYB_20__1_), .S(SUMB_20__1_) );
  AD1V2C_8TH40 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), 
        .CO(CARRYB_20__2_), .S(SUMB_20__2_) );
  AD1V2C_8TH40 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), 
        .CO(CARRYB_20__3_), .S(SUMB_20__3_) );
  AD1V2C_8TH40 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), 
        .CO(CARRYB_20__4_), .S(SUMB_20__4_) );
  AD1V2C_8TH40 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), 
        .CO(CARRYB_20__5_), .S(SUMB_20__5_) );
  AD1V2C_8TH40 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), 
        .CO(CARRYB_20__6_), .S(SUMB_20__6_) );
  AD1V2C_8TH40 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), 
        .CO(CARRYB_20__7_), .S(SUMB_20__7_) );
  AD1V2C_8TH40 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), 
        .CO(CARRYB_20__8_), .S(SUMB_20__8_) );
  AD1V2C_8TH40 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), 
        .CO(CARRYB_20__9_), .S(SUMB_20__9_) );
  AD1V2C_8TH40 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  AD1V2C_8TH40 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(CARRYB_20__11_), .S(SUMB_20__11_) );
  AD1V2C_8TH40 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(CARRYB_20__12_), .S(SUMB_20__12_) );
  AD1V2C_8TH40 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(CARRYB_20__13_), .S(SUMB_20__13_) );
  AD1V2C_8TH40 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(CARRYB_20__14_), .S(SUMB_20__14_) );
  AD1V2C_8TH40 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(CARRYB_20__15_), .S(SUMB_20__15_) );
  AD1V2C_8TH40 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(CARRYB_20__16_), .S(SUMB_20__16_) );
  AD1V2C_8TH40 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(CARRYB_20__17_), .S(SUMB_20__17_) );
  AD1V2C_8TH40 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(CARRYB_20__18_), .S(SUMB_20__18_) );
  AD1V2C_8TH40 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(CARRYB_20__19_), .S(SUMB_20__19_) );
  AD1V2C_8TH40 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(CARRYB_20__20_), .S(SUMB_20__20_) );
  AD1V2C_8TH40 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(CARRYB_20__21_), .S(SUMB_20__21_) );
  AD1V2C_8TH40 S2_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(SUMB_19__23_), .CO(CARRYB_20__22_), .S(SUMB_20__22_) );
  AD1V2C_8TH40 S2_20_23 ( .A(ab_20__23_), .B(CARRYB_19__23_), .CI(SUMB_19__24_), .CO(CARRYB_20__23_), .S(SUMB_20__23_) );
  AD1V2C_8TH40 S2_20_24 ( .A(ab_20__24_), .B(CARRYB_19__24_), .CI(SUMB_19__25_), .CO(CARRYB_20__24_), .S(SUMB_20__24_) );
  AD1V2C_8TH40 S2_20_25 ( .A(ab_20__25_), .B(CARRYB_19__25_), .CI(SUMB_19__26_), .CO(CARRYB_20__25_), .S(SUMB_20__25_) );
  AD1V2C_8TH40 S2_20_26 ( .A(ab_20__26_), .B(CARRYB_19__26_), .CI(SUMB_19__27_), .CO(CARRYB_20__26_), .S(SUMB_20__26_) );
  AD1V2C_8TH40 S2_20_27 ( .A(ab_20__27_), .B(CARRYB_19__27_), .CI(SUMB_19__28_), .CO(CARRYB_20__27_), .S(SUMB_20__27_) );
  AD1V2C_8TH40 S2_20_28 ( .A(ab_20__28_), .B(CARRYB_19__28_), .CI(SUMB_19__29_), .CO(CARRYB_20__28_), .S(SUMB_20__28_) );
  AD1V2C_8TH40 S2_20_29 ( .A(ab_20__29_), .B(CARRYB_19__29_), .CI(SUMB_19__30_), .CO(CARRYB_20__29_), .S(SUMB_20__29_) );
  AD1V2C_8TH40 S3_20_30 ( .A(ab_20__30_), .B(CARRYB_19__30_), .CI(ab_19__31_), 
        .CO(CARRYB_20__30_), .S(SUMB_20__30_) );
  AD1V2C_8TH40 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), 
        .CO(CARRYB_19__0_), .S(A1_17_) );
  AD1V2C_8TH40 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), 
        .CO(CARRYB_19__1_), .S(SUMB_19__1_) );
  AD1V2C_8TH40 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), 
        .CO(CARRYB_19__2_), .S(SUMB_19__2_) );
  AD1V2C_8TH40 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), 
        .CO(CARRYB_19__3_), .S(SUMB_19__3_) );
  AD1V2C_8TH40 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), 
        .CO(CARRYB_19__4_), .S(SUMB_19__4_) );
  AD1V2C_8TH40 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), 
        .CO(CARRYB_19__5_), .S(SUMB_19__5_) );
  AD1V2C_8TH40 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), 
        .CO(CARRYB_19__6_), .S(SUMB_19__6_) );
  AD1V2C_8TH40 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), 
        .CO(CARRYB_19__7_), .S(SUMB_19__7_) );
  AD1V2C_8TH40 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), 
        .CO(CARRYB_19__8_), .S(SUMB_19__8_) );
  AD1V2C_8TH40 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), 
        .CO(CARRYB_19__9_), .S(SUMB_19__9_) );
  AD1V2C_8TH40 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  AD1V2C_8TH40 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  AD1V2C_8TH40 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(CARRYB_19__12_), .S(SUMB_19__12_) );
  AD1V2C_8TH40 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(CARRYB_19__13_), .S(SUMB_19__13_) );
  AD1V2C_8TH40 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(CARRYB_19__14_), .S(SUMB_19__14_) );
  AD1V2C_8TH40 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(CARRYB_19__15_), .S(SUMB_19__15_) );
  AD1V2C_8TH40 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(CARRYB_19__16_), .S(SUMB_19__16_) );
  AD1V2C_8TH40 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(CARRYB_19__17_), .S(SUMB_19__17_) );
  AD1V2C_8TH40 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(CARRYB_19__18_), .S(SUMB_19__18_) );
  AD1V2C_8TH40 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(CARRYB_19__19_), .S(SUMB_19__19_) );
  AD1V2C_8TH40 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(CARRYB_19__20_), .S(SUMB_19__20_) );
  AD1V2C_8TH40 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(CARRYB_19__21_), .S(SUMB_19__21_) );
  AD1V2C_8TH40 S2_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(SUMB_18__23_), .CO(CARRYB_19__22_), .S(SUMB_19__22_) );
  AD1V2C_8TH40 S2_19_23 ( .A(ab_19__23_), .B(CARRYB_18__23_), .CI(SUMB_18__24_), .CO(CARRYB_19__23_), .S(SUMB_19__23_) );
  AD1V2C_8TH40 S2_19_24 ( .A(ab_19__24_), .B(CARRYB_18__24_), .CI(SUMB_18__25_), .CO(CARRYB_19__24_), .S(SUMB_19__24_) );
  AD1V2C_8TH40 S2_19_25 ( .A(ab_19__25_), .B(CARRYB_18__25_), .CI(SUMB_18__26_), .CO(CARRYB_19__25_), .S(SUMB_19__25_) );
  AD1V2C_8TH40 S2_19_26 ( .A(ab_19__26_), .B(CARRYB_18__26_), .CI(SUMB_18__27_), .CO(CARRYB_19__26_), .S(SUMB_19__26_) );
  AD1V2C_8TH40 S2_19_27 ( .A(ab_19__27_), .B(CARRYB_18__27_), .CI(SUMB_18__28_), .CO(CARRYB_19__27_), .S(SUMB_19__27_) );
  AD1V2C_8TH40 S2_19_28 ( .A(ab_19__28_), .B(CARRYB_18__28_), .CI(SUMB_18__29_), .CO(CARRYB_19__28_), .S(SUMB_19__28_) );
  AD1V2C_8TH40 S2_19_29 ( .A(ab_19__29_), .B(CARRYB_18__29_), .CI(SUMB_18__30_), .CO(CARRYB_19__29_), .S(SUMB_19__29_) );
  AD1V2C_8TH40 S3_19_30 ( .A(ab_19__30_), .B(CARRYB_18__30_), .CI(ab_18__31_), 
        .CO(CARRYB_19__30_), .S(SUMB_19__30_) );
  AD1V2C_8TH40 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), 
        .CO(CARRYB_18__0_), .S(A1_16_) );
  AD1V2C_8TH40 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), 
        .CO(CARRYB_18__1_), .S(SUMB_18__1_) );
  AD1V2C_8TH40 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), 
        .CO(CARRYB_18__2_), .S(SUMB_18__2_) );
  AD1V2C_8TH40 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), 
        .CO(CARRYB_18__3_), .S(SUMB_18__3_) );
  AD1V2C_8TH40 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), 
        .CO(CARRYB_18__4_), .S(SUMB_18__4_) );
  AD1V2C_8TH40 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), 
        .CO(CARRYB_18__5_), .S(SUMB_18__5_) );
  AD1V2C_8TH40 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), 
        .CO(CARRYB_18__6_), .S(SUMB_18__6_) );
  AD1V2C_8TH40 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), 
        .CO(CARRYB_18__7_), .S(SUMB_18__7_) );
  AD1V2C_8TH40 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), 
        .CO(CARRYB_18__8_), .S(SUMB_18__8_) );
  AD1V2C_8TH40 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), 
        .CO(CARRYB_18__9_), .S(SUMB_18__9_) );
  AD1V2C_8TH40 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  AD1V2C_8TH40 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  AD1V2C_8TH40 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  AD1V2C_8TH40 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(CARRYB_18__13_), .S(SUMB_18__13_) );
  AD1V2C_8TH40 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(CARRYB_18__14_), .S(SUMB_18__14_) );
  AD1V2C_8TH40 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(CARRYB_18__15_), .S(SUMB_18__15_) );
  AD1V2C_8TH40 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(CARRYB_18__16_), .S(SUMB_18__16_) );
  AD1V2C_8TH40 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(CARRYB_18__17_), .S(SUMB_18__17_) );
  AD1V2C_8TH40 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(CARRYB_18__18_), .S(SUMB_18__18_) );
  AD1V2C_8TH40 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(CARRYB_18__19_), .S(SUMB_18__19_) );
  AD1V2C_8TH40 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(CARRYB_18__20_), .S(SUMB_18__20_) );
  AD1V2C_8TH40 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(CARRYB_18__21_), .S(SUMB_18__21_) );
  AD1V2C_8TH40 S2_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(SUMB_17__23_), .CO(CARRYB_18__22_), .S(SUMB_18__22_) );
  AD1V2C_8TH40 S2_18_23 ( .A(ab_18__23_), .B(CARRYB_17__23_), .CI(SUMB_17__24_), .CO(CARRYB_18__23_), .S(SUMB_18__23_) );
  AD1V2C_8TH40 S2_18_24 ( .A(ab_18__24_), .B(CARRYB_17__24_), .CI(SUMB_17__25_), .CO(CARRYB_18__24_), .S(SUMB_18__24_) );
  AD1V2C_8TH40 S2_18_25 ( .A(ab_18__25_), .B(CARRYB_17__25_), .CI(SUMB_17__26_), .CO(CARRYB_18__25_), .S(SUMB_18__25_) );
  AD1V2C_8TH40 S2_18_26 ( .A(ab_18__26_), .B(CARRYB_17__26_), .CI(SUMB_17__27_), .CO(CARRYB_18__26_), .S(SUMB_18__26_) );
  AD1V2C_8TH40 S2_18_27 ( .A(ab_18__27_), .B(CARRYB_17__27_), .CI(SUMB_17__28_), .CO(CARRYB_18__27_), .S(SUMB_18__27_) );
  AD1V2C_8TH40 S2_18_28 ( .A(ab_18__28_), .B(CARRYB_17__28_), .CI(SUMB_17__29_), .CO(CARRYB_18__28_), .S(SUMB_18__28_) );
  AD1V2C_8TH40 S2_18_29 ( .A(ab_18__29_), .B(CARRYB_17__29_), .CI(SUMB_17__30_), .CO(CARRYB_18__29_), .S(SUMB_18__29_) );
  AD1V2C_8TH40 S3_18_30 ( .A(ab_18__30_), .B(CARRYB_17__30_), .CI(ab_17__31_), 
        .CO(CARRYB_18__30_), .S(SUMB_18__30_) );
  AD1V2C_8TH40 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), 
        .CO(CARRYB_17__0_), .S(A1_15_) );
  AD1V2C_8TH40 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), 
        .CO(CARRYB_17__1_), .S(SUMB_17__1_) );
  AD1V2C_8TH40 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), 
        .CO(CARRYB_17__2_), .S(SUMB_17__2_) );
  AD1V2C_8TH40 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), 
        .CO(CARRYB_17__3_), .S(SUMB_17__3_) );
  AD1V2C_8TH40 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), 
        .CO(CARRYB_17__4_), .S(SUMB_17__4_) );
  AD1V2C_8TH40 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), 
        .CO(CARRYB_17__5_), .S(SUMB_17__5_) );
  AD1V2C_8TH40 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), 
        .CO(CARRYB_17__6_), .S(SUMB_17__6_) );
  AD1V2C_8TH40 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), 
        .CO(CARRYB_17__7_), .S(SUMB_17__7_) );
  AD1V2C_8TH40 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), 
        .CO(CARRYB_17__8_), .S(SUMB_17__8_) );
  AD1V2C_8TH40 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), 
        .CO(CARRYB_17__9_), .S(SUMB_17__9_) );
  AD1V2C_8TH40 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  AD1V2C_8TH40 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  AD1V2C_8TH40 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  AD1V2C_8TH40 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  AD1V2C_8TH40 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(CARRYB_17__14_), .S(SUMB_17__14_) );
  AD1V2C_8TH40 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(CARRYB_17__15_), .S(SUMB_17__15_) );
  AD1V2C_8TH40 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(CARRYB_17__16_), .S(SUMB_17__16_) );
  AD1V2C_8TH40 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(CARRYB_17__17_), .S(SUMB_17__17_) );
  AD1V2C_8TH40 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(CARRYB_17__18_), .S(SUMB_17__18_) );
  AD1V2C_8TH40 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(CARRYB_17__19_), .S(SUMB_17__19_) );
  AD1V2C_8TH40 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(CARRYB_17__20_), .S(SUMB_17__20_) );
  AD1V2C_8TH40 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(CARRYB_17__21_), .S(SUMB_17__21_) );
  AD1V2C_8TH40 S2_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(SUMB_16__23_), .CO(CARRYB_17__22_), .S(SUMB_17__22_) );
  AD1V2C_8TH40 S2_17_23 ( .A(ab_17__23_), .B(CARRYB_16__23_), .CI(SUMB_16__24_), .CO(CARRYB_17__23_), .S(SUMB_17__23_) );
  AD1V2C_8TH40 S2_17_24 ( .A(ab_17__24_), .B(CARRYB_16__24_), .CI(SUMB_16__25_), .CO(CARRYB_17__24_), .S(SUMB_17__24_) );
  AD1V2C_8TH40 S2_17_25 ( .A(ab_17__25_), .B(CARRYB_16__25_), .CI(SUMB_16__26_), .CO(CARRYB_17__25_), .S(SUMB_17__25_) );
  AD1V2C_8TH40 S2_17_26 ( .A(ab_17__26_), .B(CARRYB_16__26_), .CI(SUMB_16__27_), .CO(CARRYB_17__26_), .S(SUMB_17__26_) );
  AD1V2C_8TH40 S2_17_27 ( .A(ab_17__27_), .B(CARRYB_16__27_), .CI(SUMB_16__28_), .CO(CARRYB_17__27_), .S(SUMB_17__27_) );
  AD1V2C_8TH40 S2_17_28 ( .A(ab_17__28_), .B(CARRYB_16__28_), .CI(SUMB_16__29_), .CO(CARRYB_17__28_), .S(SUMB_17__28_) );
  AD1V2C_8TH40 S2_17_29 ( .A(ab_17__29_), .B(CARRYB_16__29_), .CI(SUMB_16__30_), .CO(CARRYB_17__29_), .S(SUMB_17__29_) );
  AD1V2C_8TH40 S3_17_30 ( .A(ab_17__30_), .B(CARRYB_16__30_), .CI(ab_16__31_), 
        .CO(CARRYB_17__30_), .S(SUMB_17__30_) );
  AD1V2C_8TH40 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), 
        .CO(CARRYB_16__0_), .S(A1_14_) );
  AD1V2C_8TH40 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), 
        .CO(CARRYB_16__1_), .S(SUMB_16__1_) );
  AD1V2C_8TH40 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), 
        .CO(CARRYB_16__2_), .S(SUMB_16__2_) );
  AD1V2C_8TH40 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), 
        .CO(CARRYB_16__3_), .S(SUMB_16__3_) );
  AD1V2C_8TH40 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), 
        .CO(CARRYB_16__4_), .S(SUMB_16__4_) );
  AD1V2C_8TH40 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), 
        .CO(CARRYB_16__5_), .S(SUMB_16__5_) );
  AD1V2C_8TH40 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), 
        .CO(CARRYB_16__6_), .S(SUMB_16__6_) );
  AD1V2C_8TH40 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), 
        .CO(CARRYB_16__7_), .S(SUMB_16__7_) );
  AD1V2C_8TH40 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), 
        .CO(CARRYB_16__8_), .S(SUMB_16__8_) );
  AD1V2C_8TH40 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), 
        .CO(CARRYB_16__9_), .S(SUMB_16__9_) );
  AD1V2C_8TH40 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  AD1V2C_8TH40 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  AD1V2C_8TH40 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  AD1V2C_8TH40 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  AD1V2C_8TH40 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  AD1V2C_8TH40 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(CARRYB_16__15_), .S(SUMB_16__15_) );
  AD1V2C_8TH40 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(CARRYB_16__16_), .S(SUMB_16__16_) );
  AD1V2C_8TH40 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(CARRYB_16__17_), .S(SUMB_16__17_) );
  AD1V2C_8TH40 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(CARRYB_16__18_), .S(SUMB_16__18_) );
  AD1V2C_8TH40 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(CARRYB_16__19_), .S(SUMB_16__19_) );
  AD1V2C_8TH40 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(CARRYB_16__20_), .S(SUMB_16__20_) );
  AD1V2C_8TH40 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(CARRYB_16__21_), .S(SUMB_16__21_) );
  AD1V2C_8TH40 S2_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(SUMB_15__23_), .CO(CARRYB_16__22_), .S(SUMB_16__22_) );
  AD1V2C_8TH40 S2_16_23 ( .A(ab_16__23_), .B(CARRYB_15__23_), .CI(SUMB_15__24_), .CO(CARRYB_16__23_), .S(SUMB_16__23_) );
  AD1V2C_8TH40 S2_16_24 ( .A(ab_16__24_), .B(CARRYB_15__24_), .CI(SUMB_15__25_), .CO(CARRYB_16__24_), .S(SUMB_16__24_) );
  AD1V2C_8TH40 S2_16_25 ( .A(ab_16__25_), .B(CARRYB_15__25_), .CI(SUMB_15__26_), .CO(CARRYB_16__25_), .S(SUMB_16__25_) );
  AD1V2C_8TH40 S2_16_26 ( .A(ab_16__26_), .B(CARRYB_15__26_), .CI(SUMB_15__27_), .CO(CARRYB_16__26_), .S(SUMB_16__26_) );
  AD1V2C_8TH40 S2_16_27 ( .A(ab_16__27_), .B(CARRYB_15__27_), .CI(SUMB_15__28_), .CO(CARRYB_16__27_), .S(SUMB_16__27_) );
  AD1V2C_8TH40 S2_16_28 ( .A(ab_16__28_), .B(CARRYB_15__28_), .CI(SUMB_15__29_), .CO(CARRYB_16__28_), .S(SUMB_16__28_) );
  AD1V2C_8TH40 S2_16_29 ( .A(ab_16__29_), .B(CARRYB_15__29_), .CI(SUMB_15__30_), .CO(CARRYB_16__29_), .S(SUMB_16__29_) );
  AD1V2C_8TH40 S3_16_30 ( .A(ab_16__30_), .B(CARRYB_15__30_), .CI(ab_15__31_), 
        .CO(CARRYB_16__30_), .S(SUMB_16__30_) );
  AD1V2C_8TH40 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), 
        .CO(CARRYB_15__0_), .S(A1_13_) );
  AD1V2C_8TH40 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), 
        .CO(CARRYB_15__1_), .S(SUMB_15__1_) );
  AD1V2C_8TH40 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), 
        .CO(CARRYB_15__2_), .S(SUMB_15__2_) );
  AD1V2C_8TH40 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), 
        .CO(CARRYB_15__3_), .S(SUMB_15__3_) );
  AD1V2C_8TH40 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), 
        .CO(CARRYB_15__4_), .S(SUMB_15__4_) );
  AD1V2C_8TH40 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), 
        .CO(CARRYB_15__5_), .S(SUMB_15__5_) );
  AD1V2C_8TH40 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), 
        .CO(CARRYB_15__6_), .S(SUMB_15__6_) );
  AD1V2C_8TH40 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), 
        .CO(CARRYB_15__7_), .S(SUMB_15__7_) );
  AD1V2C_8TH40 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), 
        .CO(CARRYB_15__8_), .S(SUMB_15__8_) );
  AD1V2C_8TH40 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), 
        .CO(CARRYB_15__9_), .S(SUMB_15__9_) );
  AD1V2C_8TH40 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  AD1V2C_8TH40 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  AD1V2C_8TH40 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  AD1V2C_8TH40 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  AD1V2C_8TH40 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  AD1V2C_8TH40 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(CARRYB_15__15_), .S(SUMB_15__15_) );
  AD1V2C_8TH40 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(CARRYB_15__16_), .S(SUMB_15__16_) );
  AD1V2C_8TH40 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(CARRYB_15__17_), .S(SUMB_15__17_) );
  AD1V2C_8TH40 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(CARRYB_15__18_), .S(SUMB_15__18_) );
  AD1V2C_8TH40 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(CARRYB_15__19_), .S(SUMB_15__19_) );
  AD1V2C_8TH40 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(CARRYB_15__20_), .S(SUMB_15__20_) );
  AD1V2C_8TH40 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(CARRYB_15__21_), .S(SUMB_15__21_) );
  AD1V2C_8TH40 S2_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(SUMB_14__23_), .CO(CARRYB_15__22_), .S(SUMB_15__22_) );
  AD1V2C_8TH40 S2_15_23 ( .A(ab_15__23_), .B(CARRYB_14__23_), .CI(SUMB_14__24_), .CO(CARRYB_15__23_), .S(SUMB_15__23_) );
  AD1V2C_8TH40 S2_15_24 ( .A(ab_15__24_), .B(CARRYB_14__24_), .CI(SUMB_14__25_), .CO(CARRYB_15__24_), .S(SUMB_15__24_) );
  AD1V2C_8TH40 S2_15_25 ( .A(ab_15__25_), .B(CARRYB_14__25_), .CI(SUMB_14__26_), .CO(CARRYB_15__25_), .S(SUMB_15__25_) );
  AD1V2C_8TH40 S2_15_26 ( .A(ab_15__26_), .B(CARRYB_14__26_), .CI(SUMB_14__27_), .CO(CARRYB_15__26_), .S(SUMB_15__26_) );
  AD1V2C_8TH40 S2_15_27 ( .A(ab_15__27_), .B(CARRYB_14__27_), .CI(SUMB_14__28_), .CO(CARRYB_15__27_), .S(SUMB_15__27_) );
  AD1V2C_8TH40 S2_15_28 ( .A(ab_15__28_), .B(CARRYB_14__28_), .CI(SUMB_14__29_), .CO(CARRYB_15__28_), .S(SUMB_15__28_) );
  AD1V2C_8TH40 S2_15_29 ( .A(ab_15__29_), .B(CARRYB_14__29_), .CI(SUMB_14__30_), .CO(CARRYB_15__29_), .S(SUMB_15__29_) );
  AD1V2C_8TH40 S3_15_30 ( .A(ab_15__30_), .B(CARRYB_14__30_), .CI(ab_14__31_), 
        .CO(CARRYB_15__30_), .S(SUMB_15__30_) );
  AD1V2C_8TH40 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), 
        .CO(CARRYB_14__0_), .S(A1_12_) );
  AD1V2C_8TH40 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), 
        .CO(CARRYB_14__1_), .S(SUMB_14__1_) );
  AD1V2C_8TH40 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), 
        .CO(CARRYB_14__2_), .S(SUMB_14__2_) );
  AD1V2C_8TH40 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), 
        .CO(CARRYB_14__3_), .S(SUMB_14__3_) );
  AD1V2C_8TH40 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), 
        .CO(CARRYB_14__4_), .S(SUMB_14__4_) );
  AD1V2C_8TH40 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), 
        .CO(CARRYB_14__5_), .S(SUMB_14__5_) );
  AD1V2C_8TH40 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), 
        .CO(CARRYB_14__6_), .S(SUMB_14__6_) );
  AD1V2C_8TH40 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), 
        .CO(CARRYB_14__7_), .S(SUMB_14__7_) );
  AD1V2C_8TH40 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), 
        .CO(CARRYB_14__8_), .S(SUMB_14__8_) );
  AD1V2C_8TH40 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), 
        .CO(CARRYB_14__9_), .S(SUMB_14__9_) );
  AD1V2C_8TH40 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  AD1V2C_8TH40 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  AD1V2C_8TH40 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  AD1V2C_8TH40 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  AD1V2C_8TH40 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(CARRYB_14__14_), .S(SUMB_14__14_) );
  AD1V2C_8TH40 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  AD1V2C_8TH40 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  AD1V2C_8TH40 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(CARRYB_14__17_), .S(SUMB_14__17_) );
  AD1V2C_8TH40 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(CARRYB_14__18_), .S(SUMB_14__18_) );
  AD1V2C_8TH40 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(CARRYB_14__19_), .S(SUMB_14__19_) );
  AD1V2C_8TH40 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(CARRYB_14__20_), .S(SUMB_14__20_) );
  AD1V2C_8TH40 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(CARRYB_14__21_), .S(SUMB_14__21_) );
  AD1V2C_8TH40 S2_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(SUMB_13__23_), .CO(CARRYB_14__22_), .S(SUMB_14__22_) );
  AD1V2C_8TH40 S2_14_23 ( .A(ab_14__23_), .B(CARRYB_13__23_), .CI(SUMB_13__24_), .CO(CARRYB_14__23_), .S(SUMB_14__23_) );
  AD1V2C_8TH40 S2_14_24 ( .A(ab_14__24_), .B(CARRYB_13__24_), .CI(SUMB_13__25_), .CO(CARRYB_14__24_), .S(SUMB_14__24_) );
  AD1V2C_8TH40 S2_14_25 ( .A(ab_14__25_), .B(CARRYB_13__25_), .CI(SUMB_13__26_), .CO(CARRYB_14__25_), .S(SUMB_14__25_) );
  AD1V2C_8TH40 S2_14_26 ( .A(ab_14__26_), .B(CARRYB_13__26_), .CI(SUMB_13__27_), .CO(CARRYB_14__26_), .S(SUMB_14__26_) );
  AD1V2C_8TH40 S2_14_27 ( .A(ab_14__27_), .B(CARRYB_13__27_), .CI(SUMB_13__28_), .CO(CARRYB_14__27_), .S(SUMB_14__27_) );
  AD1V2C_8TH40 S2_14_28 ( .A(ab_14__28_), .B(CARRYB_13__28_), .CI(SUMB_13__29_), .CO(CARRYB_14__28_), .S(SUMB_14__28_) );
  AD1V2C_8TH40 S2_14_29 ( .A(ab_14__29_), .B(CARRYB_13__29_), .CI(SUMB_13__30_), .CO(CARRYB_14__29_), .S(SUMB_14__29_) );
  AD1V2C_8TH40 S3_14_30 ( .A(ab_14__30_), .B(CARRYB_13__30_), .CI(ab_13__31_), 
        .CO(CARRYB_14__30_), .S(SUMB_14__30_) );
  AD1V2C_8TH40 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), 
        .CO(CARRYB_13__0_), .S(A1_11_) );
  AD1V2C_8TH40 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), 
        .CO(CARRYB_13__1_), .S(SUMB_13__1_) );
  AD1V2C_8TH40 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), 
        .CO(CARRYB_13__2_), .S(SUMB_13__2_) );
  AD1V2C_8TH40 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), 
        .CO(CARRYB_13__3_), .S(SUMB_13__3_) );
  AD1V2C_8TH40 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), 
        .CO(CARRYB_13__4_), .S(SUMB_13__4_) );
  AD1V2C_8TH40 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), 
        .CO(CARRYB_13__5_), .S(SUMB_13__5_) );
  AD1V2C_8TH40 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), 
        .CO(CARRYB_13__6_), .S(SUMB_13__6_) );
  AD1V2C_8TH40 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), 
        .CO(CARRYB_13__7_), .S(SUMB_13__7_) );
  AD1V2C_8TH40 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), 
        .CO(CARRYB_13__8_), .S(SUMB_13__8_) );
  AD1V2C_8TH40 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), 
        .CO(CARRYB_13__9_), .S(SUMB_13__9_) );
  AD1V2C_8TH40 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  AD1V2C_8TH40 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  AD1V2C_8TH40 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  AD1V2C_8TH40 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(CARRYB_13__13_), .S(SUMB_13__13_) );
  AD1V2C_8TH40 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  AD1V2C_8TH40 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  AD1V2C_8TH40 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  AD1V2C_8TH40 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  AD1V2C_8TH40 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(CARRYB_13__18_), .S(SUMB_13__18_) );
  AD1V2C_8TH40 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(CARRYB_13__19_), .S(SUMB_13__19_) );
  AD1V2C_8TH40 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(CARRYB_13__20_), .S(SUMB_13__20_) );
  AD1V2C_8TH40 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(CARRYB_13__21_), .S(SUMB_13__21_) );
  AD1V2C_8TH40 S2_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(SUMB_12__23_), .CO(CARRYB_13__22_), .S(SUMB_13__22_) );
  AD1V2C_8TH40 S2_13_23 ( .A(ab_13__23_), .B(CARRYB_12__23_), .CI(SUMB_12__24_), .CO(CARRYB_13__23_), .S(SUMB_13__23_) );
  AD1V2C_8TH40 S2_13_24 ( .A(ab_13__24_), .B(CARRYB_12__24_), .CI(SUMB_12__25_), .CO(CARRYB_13__24_), .S(SUMB_13__24_) );
  AD1V2C_8TH40 S2_13_25 ( .A(ab_13__25_), .B(CARRYB_12__25_), .CI(SUMB_12__26_), .CO(CARRYB_13__25_), .S(SUMB_13__25_) );
  AD1V2C_8TH40 S2_13_26 ( .A(ab_13__26_), .B(CARRYB_12__26_), .CI(SUMB_12__27_), .CO(CARRYB_13__26_), .S(SUMB_13__26_) );
  AD1V2C_8TH40 S2_13_27 ( .A(ab_13__27_), .B(CARRYB_12__27_), .CI(SUMB_12__28_), .CO(CARRYB_13__27_), .S(SUMB_13__27_) );
  AD1V2C_8TH40 S2_13_28 ( .A(ab_13__28_), .B(CARRYB_12__28_), .CI(SUMB_12__29_), .CO(CARRYB_13__28_), .S(SUMB_13__28_) );
  AD1V2C_8TH40 S2_13_29 ( .A(ab_13__29_), .B(CARRYB_12__29_), .CI(SUMB_12__30_), .CO(CARRYB_13__29_), .S(SUMB_13__29_) );
  AD1V2C_8TH40 S3_13_30 ( .A(ab_13__30_), .B(CARRYB_12__30_), .CI(ab_12__31_), 
        .CO(CARRYB_13__30_), .S(SUMB_13__30_) );
  AD1V2C_8TH40 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), 
        .CO(CARRYB_12__0_), .S(A1_10_) );
  AD1V2C_8TH40 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), 
        .CO(CARRYB_12__1_), .S(SUMB_12__1_) );
  AD1V2C_8TH40 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), 
        .CO(CARRYB_12__2_), .S(SUMB_12__2_) );
  AD1V2C_8TH40 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), 
        .CO(CARRYB_12__3_), .S(SUMB_12__3_) );
  AD1V2C_8TH40 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), 
        .CO(CARRYB_12__4_), .S(SUMB_12__4_) );
  AD1V2C_8TH40 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), 
        .CO(CARRYB_12__5_), .S(SUMB_12__5_) );
  AD1V2C_8TH40 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), 
        .CO(CARRYB_12__6_), .S(SUMB_12__6_) );
  AD1V2C_8TH40 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), 
        .CO(CARRYB_12__7_), .S(SUMB_12__7_) );
  AD1V2C_8TH40 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), 
        .CO(CARRYB_12__8_), .S(SUMB_12__8_) );
  AD1V2C_8TH40 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), 
        .CO(CARRYB_12__9_), .S(SUMB_12__9_) );
  AD1V2C_8TH40 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  AD1V2C_8TH40 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  AD1V2C_8TH40 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(CARRYB_12__12_), .S(SUMB_12__12_) );
  AD1V2C_8TH40 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  AD1V2C_8TH40 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  AD1V2C_8TH40 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  AD1V2C_8TH40 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  AD1V2C_8TH40 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  AD1V2C_8TH40 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  AD1V2C_8TH40 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(CARRYB_12__19_), .S(SUMB_12__19_) );
  AD1V2C_8TH40 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(CARRYB_12__20_), .S(SUMB_12__20_) );
  AD1V2C_8TH40 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(CARRYB_12__21_), .S(SUMB_12__21_) );
  AD1V2C_8TH40 S2_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(SUMB_11__23_), .CO(CARRYB_12__22_), .S(SUMB_12__22_) );
  AD1V2C_8TH40 S2_12_23 ( .A(ab_12__23_), .B(CARRYB_11__23_), .CI(SUMB_11__24_), .CO(CARRYB_12__23_), .S(SUMB_12__23_) );
  AD1V2C_8TH40 S2_12_24 ( .A(ab_12__24_), .B(CARRYB_11__24_), .CI(SUMB_11__25_), .CO(CARRYB_12__24_), .S(SUMB_12__24_) );
  AD1V2C_8TH40 S2_12_25 ( .A(ab_12__25_), .B(CARRYB_11__25_), .CI(SUMB_11__26_), .CO(CARRYB_12__25_), .S(SUMB_12__25_) );
  AD1V2C_8TH40 S2_12_26 ( .A(ab_12__26_), .B(CARRYB_11__26_), .CI(SUMB_11__27_), .CO(CARRYB_12__26_), .S(SUMB_12__26_) );
  AD1V2C_8TH40 S2_12_27 ( .A(ab_12__27_), .B(CARRYB_11__27_), .CI(SUMB_11__28_), .CO(CARRYB_12__27_), .S(SUMB_12__27_) );
  AD1V2C_8TH40 S2_12_28 ( .A(ab_12__28_), .B(CARRYB_11__28_), .CI(SUMB_11__29_), .CO(CARRYB_12__28_), .S(SUMB_12__28_) );
  AD1V2C_8TH40 S2_12_29 ( .A(ab_12__29_), .B(CARRYB_11__29_), .CI(SUMB_11__30_), .CO(CARRYB_12__29_), .S(SUMB_12__29_) );
  AD1V2C_8TH40 S3_12_30 ( .A(ab_12__30_), .B(CARRYB_11__30_), .CI(ab_11__31_), 
        .CO(CARRYB_12__30_), .S(SUMB_12__30_) );
  AD1V2C_8TH40 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), 
        .CO(CARRYB_11__0_), .S(A1_9_) );
  AD1V2C_8TH40 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), 
        .CO(CARRYB_11__1_), .S(SUMB_11__1_) );
  AD1V2C_8TH40 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), 
        .CO(CARRYB_11__2_), .S(SUMB_11__2_) );
  AD1V2C_8TH40 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), 
        .CO(CARRYB_11__3_), .S(SUMB_11__3_) );
  AD1V2C_8TH40 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), 
        .CO(CARRYB_11__4_), .S(SUMB_11__4_) );
  AD1V2C_8TH40 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), 
        .CO(CARRYB_11__5_), .S(SUMB_11__5_) );
  AD1V2C_8TH40 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), 
        .CO(CARRYB_11__6_), .S(SUMB_11__6_) );
  AD1V2C_8TH40 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), 
        .CO(CARRYB_11__7_), .S(SUMB_11__7_) );
  AD1V2C_8TH40 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), 
        .CO(CARRYB_11__8_), .S(SUMB_11__8_) );
  AD1V2C_8TH40 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), 
        .CO(CARRYB_11__9_), .S(SUMB_11__9_) );
  AD1V2C_8TH40 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  AD1V2C_8TH40 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(CARRYB_11__11_), .S(SUMB_11__11_) );
  AD1V2C_8TH40 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  AD1V2C_8TH40 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  AD1V2C_8TH40 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  AD1V2C_8TH40 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  AD1V2C_8TH40 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  AD1V2C_8TH40 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  AD1V2C_8TH40 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  AD1V2C_8TH40 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  AD1V2C_8TH40 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(CARRYB_11__20_), .S(SUMB_11__20_) );
  AD1V2C_8TH40 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(CARRYB_11__21_), .S(SUMB_11__21_) );
  AD1V2C_8TH40 S2_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(SUMB_10__23_), .CO(CARRYB_11__22_), .S(SUMB_11__22_) );
  AD1V2C_8TH40 S2_11_23 ( .A(ab_11__23_), .B(CARRYB_10__23_), .CI(SUMB_10__24_), .CO(CARRYB_11__23_), .S(SUMB_11__23_) );
  AD1V2C_8TH40 S2_11_24 ( .A(ab_11__24_), .B(CARRYB_10__24_), .CI(SUMB_10__25_), .CO(CARRYB_11__24_), .S(SUMB_11__24_) );
  AD1V2C_8TH40 S2_11_25 ( .A(ab_11__25_), .B(CARRYB_10__25_), .CI(SUMB_10__26_), .CO(CARRYB_11__25_), .S(SUMB_11__25_) );
  AD1V2C_8TH40 S2_11_26 ( .A(ab_11__26_), .B(CARRYB_10__26_), .CI(SUMB_10__27_), .CO(CARRYB_11__26_), .S(SUMB_11__26_) );
  AD1V2C_8TH40 S2_11_27 ( .A(ab_11__27_), .B(CARRYB_10__27_), .CI(SUMB_10__28_), .CO(CARRYB_11__27_), .S(SUMB_11__27_) );
  AD1V2C_8TH40 S2_11_28 ( .A(ab_11__28_), .B(CARRYB_10__28_), .CI(SUMB_10__29_), .CO(CARRYB_11__28_), .S(SUMB_11__28_) );
  AD1V2C_8TH40 S2_11_29 ( .A(ab_11__29_), .B(CARRYB_10__29_), .CI(SUMB_10__30_), .CO(CARRYB_11__29_), .S(SUMB_11__29_) );
  AD1V2C_8TH40 S3_11_30 ( .A(ab_11__30_), .B(CARRYB_10__30_), .CI(ab_10__31_), 
        .CO(CARRYB_11__30_), .S(SUMB_11__30_) );
  AD1V2C_8TH40 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), 
        .CO(CARRYB_10__0_), .S(A1_8_) );
  AD1V2C_8TH40 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), 
        .CO(CARRYB_10__1_), .S(SUMB_10__1_) );
  AD1V2C_8TH40 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), 
        .CO(CARRYB_10__2_), .S(SUMB_10__2_) );
  AD1V2C_8TH40 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), 
        .CO(CARRYB_10__3_), .S(SUMB_10__3_) );
  AD1V2C_8TH40 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), 
        .CO(CARRYB_10__4_), .S(SUMB_10__4_) );
  AD1V2C_8TH40 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), 
        .CO(CARRYB_10__5_), .S(SUMB_10__5_) );
  AD1V2C_8TH40 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), 
        .CO(CARRYB_10__6_), .S(SUMB_10__6_) );
  AD1V2C_8TH40 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), 
        .CO(CARRYB_10__7_), .S(SUMB_10__7_) );
  AD1V2C_8TH40 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), 
        .CO(CARRYB_10__8_), .S(SUMB_10__8_) );
  AD1V2C_8TH40 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), 
        .CO(CARRYB_10__9_), .S(SUMB_10__9_) );
  AD1V2C_8TH40 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), 
        .CO(CARRYB_10__10_), .S(SUMB_10__10_) );
  AD1V2C_8TH40 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), 
        .CO(CARRYB_10__11_), .S(SUMB_10__11_) );
  AD1V2C_8TH40 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), 
        .CO(CARRYB_10__12_), .S(SUMB_10__12_) );
  AD1V2C_8TH40 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), 
        .CO(CARRYB_10__13_), .S(SUMB_10__13_) );
  AD1V2C_8TH40 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), 
        .CO(CARRYB_10__14_), .S(SUMB_10__14_) );
  AD1V2C_8TH40 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), 
        .CO(CARRYB_10__15_), .S(SUMB_10__15_) );
  AD1V2C_8TH40 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), 
        .CO(CARRYB_10__16_), .S(SUMB_10__16_) );
  AD1V2C_8TH40 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), 
        .CO(CARRYB_10__17_), .S(SUMB_10__17_) );
  AD1V2C_8TH40 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), 
        .CO(CARRYB_10__18_), .S(SUMB_10__18_) );
  AD1V2C_8TH40 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), 
        .CO(CARRYB_10__19_), .S(SUMB_10__19_) );
  AD1V2C_8TH40 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), 
        .CO(CARRYB_10__20_), .S(SUMB_10__20_) );
  AD1V2C_8TH40 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), 
        .CO(CARRYB_10__21_), .S(SUMB_10__21_) );
  AD1V2C_8TH40 S2_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(SUMB_9__23_), 
        .CO(CARRYB_10__22_), .S(SUMB_10__22_) );
  AD1V2C_8TH40 S2_10_23 ( .A(ab_10__23_), .B(CARRYB_9__23_), .CI(SUMB_9__24_), 
        .CO(CARRYB_10__23_), .S(SUMB_10__23_) );
  AD1V2C_8TH40 S2_10_24 ( .A(ab_10__24_), .B(CARRYB_9__24_), .CI(SUMB_9__25_), 
        .CO(CARRYB_10__24_), .S(SUMB_10__24_) );
  AD1V2C_8TH40 S2_10_25 ( .A(ab_10__25_), .B(CARRYB_9__25_), .CI(SUMB_9__26_), 
        .CO(CARRYB_10__25_), .S(SUMB_10__25_) );
  AD1V2C_8TH40 S2_10_26 ( .A(ab_10__26_), .B(CARRYB_9__26_), .CI(SUMB_9__27_), 
        .CO(CARRYB_10__26_), .S(SUMB_10__26_) );
  AD1V2C_8TH40 S2_10_27 ( .A(ab_10__27_), .B(CARRYB_9__27_), .CI(SUMB_9__28_), 
        .CO(CARRYB_10__27_), .S(SUMB_10__27_) );
  AD1V2C_8TH40 S2_10_28 ( .A(ab_10__28_), .B(CARRYB_9__28_), .CI(SUMB_9__29_), 
        .CO(CARRYB_10__28_), .S(SUMB_10__28_) );
  AD1V2C_8TH40 S2_10_29 ( .A(ab_10__29_), .B(CARRYB_9__29_), .CI(SUMB_9__30_), 
        .CO(CARRYB_10__29_), .S(SUMB_10__29_) );
  AD1V2C_8TH40 S3_10_30 ( .A(ab_10__30_), .B(CARRYB_9__30_), .CI(ab_9__31_), 
        .CO(CARRYB_10__30_), .S(SUMB_10__30_) );
  AD1V2C_8TH40 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  AD1V2C_8TH40 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  AD1V2C_8TH40 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  AD1V2C_8TH40 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  AD1V2C_8TH40 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  AD1V2C_8TH40 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  AD1V2C_8TH40 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  AD1V2C_8TH40 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  AD1V2C_8TH40 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  AD1V2C_8TH40 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  AD1V2C_8TH40 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), 
        .CO(CARRYB_9__10_), .S(SUMB_9__10_) );
  AD1V2C_8TH40 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), 
        .CO(CARRYB_9__11_), .S(SUMB_9__11_) );
  AD1V2C_8TH40 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), 
        .CO(CARRYB_9__12_), .S(SUMB_9__12_) );
  AD1V2C_8TH40 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), 
        .CO(CARRYB_9__13_), .S(SUMB_9__13_) );
  AD1V2C_8TH40 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), 
        .CO(CARRYB_9__14_), .S(SUMB_9__14_) );
  AD1V2C_8TH40 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), 
        .CO(CARRYB_9__15_), .S(SUMB_9__15_) );
  AD1V2C_8TH40 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), 
        .CO(CARRYB_9__16_), .S(SUMB_9__16_) );
  AD1V2C_8TH40 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), 
        .CO(CARRYB_9__17_), .S(SUMB_9__17_) );
  AD1V2C_8TH40 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), 
        .CO(CARRYB_9__18_), .S(SUMB_9__18_) );
  AD1V2C_8TH40 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), 
        .CO(CARRYB_9__19_), .S(SUMB_9__19_) );
  AD1V2C_8TH40 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), 
        .CO(CARRYB_9__20_), .S(SUMB_9__20_) );
  AD1V2C_8TH40 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), 
        .CO(CARRYB_9__21_), .S(SUMB_9__21_) );
  AD1V2C_8TH40 S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), 
        .CO(CARRYB_9__22_), .S(SUMB_9__22_) );
  AD1V2C_8TH40 S2_9_23 ( .A(ab_9__23_), .B(CARRYB_8__23_), .CI(SUMB_8__24_), 
        .CO(CARRYB_9__23_), .S(SUMB_9__23_) );
  AD1V2C_8TH40 S2_9_24 ( .A(ab_9__24_), .B(CARRYB_8__24_), .CI(SUMB_8__25_), 
        .CO(CARRYB_9__24_), .S(SUMB_9__24_) );
  AD1V2C_8TH40 S2_9_25 ( .A(ab_9__25_), .B(CARRYB_8__25_), .CI(SUMB_8__26_), 
        .CO(CARRYB_9__25_), .S(SUMB_9__25_) );
  AD1V2C_8TH40 S2_9_26 ( .A(ab_9__26_), .B(CARRYB_8__26_), .CI(SUMB_8__27_), 
        .CO(CARRYB_9__26_), .S(SUMB_9__26_) );
  AD1V2C_8TH40 S2_9_27 ( .A(ab_9__27_), .B(CARRYB_8__27_), .CI(SUMB_8__28_), 
        .CO(CARRYB_9__27_), .S(SUMB_9__27_) );
  AD1V2C_8TH40 S2_9_28 ( .A(ab_9__28_), .B(CARRYB_8__28_), .CI(SUMB_8__29_), 
        .CO(CARRYB_9__28_), .S(SUMB_9__28_) );
  AD1V2C_8TH40 S2_9_29 ( .A(ab_9__29_), .B(CARRYB_8__29_), .CI(SUMB_8__30_), 
        .CO(CARRYB_9__29_), .S(SUMB_9__29_) );
  AD1V2C_8TH40 S3_9_30 ( .A(ab_9__30_), .B(CARRYB_8__30_), .CI(ab_8__31_), 
        .CO(CARRYB_9__30_), .S(SUMB_9__30_) );
  AD1V2C_8TH40 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  AD1V2C_8TH40 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  AD1V2C_8TH40 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  AD1V2C_8TH40 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  AD1V2C_8TH40 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  AD1V2C_8TH40 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  AD1V2C_8TH40 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  AD1V2C_8TH40 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  AD1V2C_8TH40 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  AD1V2C_8TH40 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  AD1V2C_8TH40 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), 
        .CO(CARRYB_8__10_), .S(SUMB_8__10_) );
  AD1V2C_8TH40 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), 
        .CO(CARRYB_8__11_), .S(SUMB_8__11_) );
  AD1V2C_8TH40 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), 
        .CO(CARRYB_8__12_), .S(SUMB_8__12_) );
  AD1V2C_8TH40 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), 
        .CO(CARRYB_8__13_), .S(SUMB_8__13_) );
  AD1V2C_8TH40 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), 
        .CO(CARRYB_8__14_), .S(SUMB_8__14_) );
  AD1V2C_8TH40 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), 
        .CO(CARRYB_8__15_), .S(SUMB_8__15_) );
  AD1V2C_8TH40 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), 
        .CO(CARRYB_8__16_), .S(SUMB_8__16_) );
  AD1V2C_8TH40 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), 
        .CO(CARRYB_8__17_), .S(SUMB_8__17_) );
  AD1V2C_8TH40 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), 
        .CO(CARRYB_8__18_), .S(SUMB_8__18_) );
  AD1V2C_8TH40 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), 
        .CO(CARRYB_8__19_), .S(SUMB_8__19_) );
  AD1V2C_8TH40 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), 
        .CO(CARRYB_8__20_), .S(SUMB_8__20_) );
  AD1V2C_8TH40 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), 
        .CO(CARRYB_8__21_), .S(SUMB_8__21_) );
  AD1V2C_8TH40 S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), 
        .CO(CARRYB_8__22_), .S(SUMB_8__22_) );
  AD1V2C_8TH40 S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), 
        .CO(CARRYB_8__23_), .S(SUMB_8__23_) );
  AD1V2C_8TH40 S2_8_24 ( .A(ab_8__24_), .B(CARRYB_7__24_), .CI(SUMB_7__25_), 
        .CO(CARRYB_8__24_), .S(SUMB_8__24_) );
  AD1V2C_8TH40 S2_8_25 ( .A(ab_8__25_), .B(CARRYB_7__25_), .CI(SUMB_7__26_), 
        .CO(CARRYB_8__25_), .S(SUMB_8__25_) );
  AD1V2C_8TH40 S2_8_26 ( .A(ab_8__26_), .B(CARRYB_7__26_), .CI(SUMB_7__27_), 
        .CO(CARRYB_8__26_), .S(SUMB_8__26_) );
  AD1V2C_8TH40 S2_8_27 ( .A(ab_8__27_), .B(CARRYB_7__27_), .CI(SUMB_7__28_), 
        .CO(CARRYB_8__27_), .S(SUMB_8__27_) );
  AD1V2C_8TH40 S2_8_28 ( .A(ab_8__28_), .B(CARRYB_7__28_), .CI(SUMB_7__29_), 
        .CO(CARRYB_8__28_), .S(SUMB_8__28_) );
  AD1V2C_8TH40 S2_8_29 ( .A(ab_8__29_), .B(CARRYB_7__29_), .CI(SUMB_7__30_), 
        .CO(CARRYB_8__29_), .S(SUMB_8__29_) );
  AD1V2C_8TH40 S3_8_30 ( .A(ab_8__30_), .B(CARRYB_7__30_), .CI(ab_7__31_), 
        .CO(CARRYB_8__30_), .S(SUMB_8__30_) );
  AD1V2C_8TH40 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  AD1V2C_8TH40 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  AD1V2C_8TH40 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  AD1V2C_8TH40 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  AD1V2C_8TH40 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  AD1V2C_8TH40 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  AD1V2C_8TH40 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  AD1V2C_8TH40 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  AD1V2C_8TH40 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  AD1V2C_8TH40 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  AD1V2C_8TH40 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), 
        .CO(CARRYB_7__10_), .S(SUMB_7__10_) );
  AD1V2C_8TH40 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), 
        .CO(CARRYB_7__11_), .S(SUMB_7__11_) );
  AD1V2C_8TH40 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), 
        .CO(CARRYB_7__12_), .S(SUMB_7__12_) );
  AD1V2C_8TH40 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), 
        .CO(CARRYB_7__13_), .S(SUMB_7__13_) );
  AD1V2C_8TH40 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), 
        .CO(CARRYB_7__14_), .S(SUMB_7__14_) );
  AD1V2C_8TH40 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), 
        .CO(CARRYB_7__15_), .S(SUMB_7__15_) );
  AD1V2C_8TH40 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), 
        .CO(CARRYB_7__16_), .S(SUMB_7__16_) );
  AD1V2C_8TH40 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), 
        .CO(CARRYB_7__17_), .S(SUMB_7__17_) );
  AD1V2C_8TH40 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), 
        .CO(CARRYB_7__18_), .S(SUMB_7__18_) );
  AD1V2C_8TH40 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), 
        .CO(CARRYB_7__19_), .S(SUMB_7__19_) );
  AD1V2C_8TH40 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), 
        .CO(CARRYB_7__20_), .S(SUMB_7__20_) );
  AD1V2C_8TH40 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), 
        .CO(CARRYB_7__21_), .S(SUMB_7__21_) );
  AD1V2C_8TH40 S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), 
        .CO(CARRYB_7__22_), .S(SUMB_7__22_) );
  AD1V2C_8TH40 S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), 
        .CO(CARRYB_7__23_), .S(SUMB_7__23_) );
  AD1V2C_8TH40 S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), 
        .CO(CARRYB_7__24_), .S(SUMB_7__24_) );
  AD1V2C_8TH40 S2_7_25 ( .A(ab_7__25_), .B(CARRYB_6__25_), .CI(SUMB_6__26_), 
        .CO(CARRYB_7__25_), .S(SUMB_7__25_) );
  AD1V2C_8TH40 S2_7_26 ( .A(ab_7__26_), .B(CARRYB_6__26_), .CI(SUMB_6__27_), 
        .CO(CARRYB_7__26_), .S(SUMB_7__26_) );
  AD1V2C_8TH40 S2_7_27 ( .A(ab_7__27_), .B(CARRYB_6__27_), .CI(SUMB_6__28_), 
        .CO(CARRYB_7__27_), .S(SUMB_7__27_) );
  AD1V2C_8TH40 S2_7_28 ( .A(ab_7__28_), .B(CARRYB_6__28_), .CI(SUMB_6__29_), 
        .CO(CARRYB_7__28_), .S(SUMB_7__28_) );
  AD1V2C_8TH40 S2_7_29 ( .A(ab_7__29_), .B(CARRYB_6__29_), .CI(SUMB_6__30_), 
        .CO(CARRYB_7__29_), .S(SUMB_7__29_) );
  AD1V2C_8TH40 S3_7_30 ( .A(ab_7__30_), .B(CARRYB_6__30_), .CI(ab_6__31_), 
        .CO(CARRYB_7__30_), .S(SUMB_7__30_) );
  AD1V2C_8TH40 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  AD1V2C_8TH40 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  AD1V2C_8TH40 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  AD1V2C_8TH40 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  AD1V2C_8TH40 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  AD1V2C_8TH40 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  AD1V2C_8TH40 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  AD1V2C_8TH40 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  AD1V2C_8TH40 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  AD1V2C_8TH40 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  AD1V2C_8TH40 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), 
        .CO(CARRYB_6__10_), .S(SUMB_6__10_) );
  AD1V2C_8TH40 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), 
        .CO(CARRYB_6__11_), .S(SUMB_6__11_) );
  AD1V2C_8TH40 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), 
        .CO(CARRYB_6__12_), .S(SUMB_6__12_) );
  AD1V2C_8TH40 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), 
        .CO(CARRYB_6__13_), .S(SUMB_6__13_) );
  AD1V2C_8TH40 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), 
        .CO(CARRYB_6__14_), .S(SUMB_6__14_) );
  AD1V2C_8TH40 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), 
        .CO(CARRYB_6__15_), .S(SUMB_6__15_) );
  AD1V2C_8TH40 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), 
        .CO(CARRYB_6__16_), .S(SUMB_6__16_) );
  AD1V2C_8TH40 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), 
        .CO(CARRYB_6__17_), .S(SUMB_6__17_) );
  AD1V2C_8TH40 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), 
        .CO(CARRYB_6__18_), .S(SUMB_6__18_) );
  AD1V2C_8TH40 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), 
        .CO(CARRYB_6__19_), .S(SUMB_6__19_) );
  AD1V2C_8TH40 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), 
        .CO(CARRYB_6__20_), .S(SUMB_6__20_) );
  AD1V2C_8TH40 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), 
        .CO(CARRYB_6__21_), .S(SUMB_6__21_) );
  AD1V2C_8TH40 S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), 
        .CO(CARRYB_6__22_), .S(SUMB_6__22_) );
  AD1V2C_8TH40 S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), 
        .CO(CARRYB_6__23_), .S(SUMB_6__23_) );
  AD1V2C_8TH40 S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), 
        .CO(CARRYB_6__24_), .S(SUMB_6__24_) );
  AD1V2C_8TH40 S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), 
        .CO(CARRYB_6__25_), .S(SUMB_6__25_) );
  AD1V2C_8TH40 S2_6_26 ( .A(ab_6__26_), .B(CARRYB_5__26_), .CI(SUMB_5__27_), 
        .CO(CARRYB_6__26_), .S(SUMB_6__26_) );
  AD1V2C_8TH40 S2_6_27 ( .A(ab_6__27_), .B(CARRYB_5__27_), .CI(SUMB_5__28_), 
        .CO(CARRYB_6__27_), .S(SUMB_6__27_) );
  AD1V2C_8TH40 S2_6_28 ( .A(ab_6__28_), .B(CARRYB_5__28_), .CI(SUMB_5__29_), 
        .CO(CARRYB_6__28_), .S(SUMB_6__28_) );
  AD1V2C_8TH40 S2_6_29 ( .A(ab_6__29_), .B(CARRYB_5__29_), .CI(SUMB_5__30_), 
        .CO(CARRYB_6__29_), .S(SUMB_6__29_) );
  AD1V2C_8TH40 S3_6_30 ( .A(ab_6__30_), .B(CARRYB_5__30_), .CI(ab_5__31_), 
        .CO(CARRYB_6__30_), .S(SUMB_6__30_) );
  AD1V2C_8TH40 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  AD1V2C_8TH40 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  AD1V2C_8TH40 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  AD1V2C_8TH40 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  AD1V2C_8TH40 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  AD1V2C_8TH40 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  AD1V2C_8TH40 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  AD1V2C_8TH40 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  AD1V2C_8TH40 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  AD1V2C_8TH40 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  AD1V2C_8TH40 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), 
        .CO(CARRYB_5__10_), .S(SUMB_5__10_) );
  AD1V2C_8TH40 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), 
        .CO(CARRYB_5__11_), .S(SUMB_5__11_) );
  AD1V2C_8TH40 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), 
        .CO(CARRYB_5__12_), .S(SUMB_5__12_) );
  AD1V2C_8TH40 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), 
        .CO(CARRYB_5__13_), .S(SUMB_5__13_) );
  AD1V2C_8TH40 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), 
        .CO(CARRYB_5__14_), .S(SUMB_5__14_) );
  AD1V2C_8TH40 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), 
        .CO(CARRYB_5__15_), .S(SUMB_5__15_) );
  AD1V2C_8TH40 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), 
        .CO(CARRYB_5__16_), .S(SUMB_5__16_) );
  AD1V2C_8TH40 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), 
        .CO(CARRYB_5__17_), .S(SUMB_5__17_) );
  AD1V2C_8TH40 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), 
        .CO(CARRYB_5__18_), .S(SUMB_5__18_) );
  AD1V2C_8TH40 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), 
        .CO(CARRYB_5__19_), .S(SUMB_5__19_) );
  AD1V2C_8TH40 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), 
        .CO(CARRYB_5__20_), .S(SUMB_5__20_) );
  AD1V2C_8TH40 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), 
        .CO(CARRYB_5__21_), .S(SUMB_5__21_) );
  AD1V2C_8TH40 S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), 
        .CO(CARRYB_5__22_), .S(SUMB_5__22_) );
  AD1V2C_8TH40 S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), 
        .CO(CARRYB_5__23_), .S(SUMB_5__23_) );
  AD1V2C_8TH40 S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), 
        .CO(CARRYB_5__24_), .S(SUMB_5__24_) );
  AD1V2C_8TH40 S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), 
        .CO(CARRYB_5__25_), .S(SUMB_5__25_) );
  AD1V2C_8TH40 S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), 
        .CO(CARRYB_5__26_), .S(SUMB_5__26_) );
  AD1V2C_8TH40 S2_5_27 ( .A(ab_5__27_), .B(CARRYB_4__27_), .CI(SUMB_4__28_), 
        .CO(CARRYB_5__27_), .S(SUMB_5__27_) );
  AD1V2C_8TH40 S2_5_28 ( .A(ab_5__28_), .B(CARRYB_4__28_), .CI(SUMB_4__29_), 
        .CO(CARRYB_5__28_), .S(SUMB_5__28_) );
  AD1V2C_8TH40 S2_5_29 ( .A(ab_5__29_), .B(CARRYB_4__29_), .CI(SUMB_4__30_), 
        .CO(CARRYB_5__29_), .S(SUMB_5__29_) );
  AD1V2C_8TH40 S3_5_30 ( .A(ab_5__30_), .B(CARRYB_4__30_), .CI(ab_4__31_), 
        .CO(CARRYB_5__30_), .S(SUMB_5__30_) );
  AD1V2C_8TH40 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  AD1V2C_8TH40 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  AD1V2C_8TH40 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  AD1V2C_8TH40 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  AD1V2C_8TH40 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  AD1V2C_8TH40 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  AD1V2C_8TH40 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  AD1V2C_8TH40 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  AD1V2C_8TH40 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  AD1V2C_8TH40 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  AD1V2C_8TH40 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), 
        .CO(CARRYB_4__10_), .S(SUMB_4__10_) );
  AD1V2C_8TH40 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), 
        .CO(CARRYB_4__11_), .S(SUMB_4__11_) );
  AD1V2C_8TH40 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), 
        .CO(CARRYB_4__12_), .S(SUMB_4__12_) );
  AD1V2C_8TH40 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), 
        .CO(CARRYB_4__13_), .S(SUMB_4__13_) );
  AD1V2C_8TH40 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), 
        .CO(CARRYB_4__14_), .S(SUMB_4__14_) );
  AD1V2C_8TH40 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), 
        .CO(CARRYB_4__15_), .S(SUMB_4__15_) );
  AD1V2C_8TH40 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), 
        .CO(CARRYB_4__16_), .S(SUMB_4__16_) );
  AD1V2C_8TH40 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), 
        .CO(CARRYB_4__17_), .S(SUMB_4__17_) );
  AD1V2C_8TH40 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), 
        .CO(CARRYB_4__18_), .S(SUMB_4__18_) );
  AD1V2C_8TH40 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), 
        .CO(CARRYB_4__19_), .S(SUMB_4__19_) );
  AD1V2C_8TH40 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), 
        .CO(CARRYB_4__20_), .S(SUMB_4__20_) );
  AD1V2C_8TH40 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), 
        .CO(CARRYB_4__21_), .S(SUMB_4__21_) );
  AD1V2C_8TH40 S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), 
        .CO(CARRYB_4__22_), .S(SUMB_4__22_) );
  AD1V2C_8TH40 S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), 
        .CO(CARRYB_4__23_), .S(SUMB_4__23_) );
  AD1V2C_8TH40 S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), 
        .CO(CARRYB_4__24_), .S(SUMB_4__24_) );
  AD1V2C_8TH40 S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), 
        .CO(CARRYB_4__25_), .S(SUMB_4__25_) );
  AD1V2C_8TH40 S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), 
        .CO(CARRYB_4__26_), .S(SUMB_4__26_) );
  AD1V2C_8TH40 S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), 
        .CO(CARRYB_4__27_), .S(SUMB_4__27_) );
  AD1V2C_8TH40 S2_4_28 ( .A(ab_4__28_), .B(CARRYB_3__28_), .CI(SUMB_3__29_), 
        .CO(CARRYB_4__28_), .S(SUMB_4__28_) );
  AD1V2C_8TH40 S2_4_29 ( .A(ab_4__29_), .B(CARRYB_3__29_), .CI(SUMB_3__30_), 
        .CO(CARRYB_4__29_), .S(SUMB_4__29_) );
  AD1V2C_8TH40 S3_4_30 ( .A(ab_4__30_), .B(CARRYB_3__30_), .CI(ab_3__31_), 
        .CO(CARRYB_4__30_), .S(SUMB_4__30_) );
  AD1V2C_8TH40 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  AD1V2C_8TH40 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  AD1V2C_8TH40 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  AD1V2C_8TH40 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  AD1V2C_8TH40 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  AD1V2C_8TH40 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  AD1V2C_8TH40 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  AD1V2C_8TH40 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  AD1V2C_8TH40 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  AD1V2C_8TH40 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  AD1V2C_8TH40 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), 
        .CO(CARRYB_3__10_), .S(SUMB_3__10_) );
  AD1V2C_8TH40 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), 
        .CO(CARRYB_3__11_), .S(SUMB_3__11_) );
  AD1V2C_8TH40 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), 
        .CO(CARRYB_3__12_), .S(SUMB_3__12_) );
  AD1V2C_8TH40 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), 
        .CO(CARRYB_3__13_), .S(SUMB_3__13_) );
  AD1V2C_8TH40 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), 
        .CO(CARRYB_3__14_), .S(SUMB_3__14_) );
  AD1V2C_8TH40 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), 
        .CO(CARRYB_3__15_), .S(SUMB_3__15_) );
  AD1V2C_8TH40 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), 
        .CO(CARRYB_3__16_), .S(SUMB_3__16_) );
  AD1V2C_8TH40 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), 
        .CO(CARRYB_3__17_), .S(SUMB_3__17_) );
  AD1V2C_8TH40 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), 
        .CO(CARRYB_3__18_), .S(SUMB_3__18_) );
  AD1V2C_8TH40 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), 
        .CO(CARRYB_3__19_), .S(SUMB_3__19_) );
  AD1V2C_8TH40 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), 
        .CO(CARRYB_3__20_), .S(SUMB_3__20_) );
  AD1V2C_8TH40 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), 
        .CO(CARRYB_3__21_), .S(SUMB_3__21_) );
  AD1V2C_8TH40 S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), 
        .CO(CARRYB_3__22_), .S(SUMB_3__22_) );
  AD1V2C_8TH40 S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), 
        .CO(CARRYB_3__23_), .S(SUMB_3__23_) );
  AD1V2C_8TH40 S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), 
        .CO(CARRYB_3__24_), .S(SUMB_3__24_) );
  AD1V2C_8TH40 S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), 
        .CO(CARRYB_3__25_), .S(SUMB_3__25_) );
  AD1V2C_8TH40 S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), 
        .CO(CARRYB_3__26_), .S(SUMB_3__26_) );
  AD1V2C_8TH40 S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), 
        .CO(CARRYB_3__27_), .S(SUMB_3__27_) );
  AD1V2C_8TH40 S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), 
        .CO(CARRYB_3__28_), .S(SUMB_3__28_) );
  AD1V2C_8TH40 S2_3_29 ( .A(ab_3__29_), .B(CARRYB_2__29_), .CI(SUMB_2__30_), 
        .CO(CARRYB_3__29_), .S(SUMB_3__29_) );
  AD1V2C_8TH40 S3_3_30 ( .A(ab_3__30_), .B(CARRYB_2__30_), .CI(ab_2__31_), 
        .CO(CARRYB_3__30_), .S(SUMB_3__30_) );
  AD1V2C_8TH40 S1_2_0 ( .A(ab_2__0_), .B(n32), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  AD1V2C_8TH40 S2_2_1 ( .A(ab_2__1_), .B(n31), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  AD1V2C_8TH40 S2_2_2 ( .A(ab_2__2_), .B(n30), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  AD1V2C_8TH40 S2_2_3 ( .A(ab_2__3_), .B(n29), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  AD1V2C_8TH40 S2_2_4 ( .A(ab_2__4_), .B(n28), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  AD1V2C_8TH40 S2_2_5 ( .A(ab_2__5_), .B(n27), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  AD1V2C_8TH40 S2_2_6 ( .A(ab_2__6_), .B(n26), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  AD1V2C_8TH40 S2_2_7 ( .A(ab_2__7_), .B(n25), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  AD1V2C_8TH40 S2_2_8 ( .A(ab_2__8_), .B(n24), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  AD1V2C_8TH40 S2_2_9 ( .A(ab_2__9_), .B(n23), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  AD1V2C_8TH40 S2_2_10 ( .A(ab_2__10_), .B(n22), .CI(SUMB_1__11_), .CO(
        CARRYB_2__10_), .S(SUMB_2__10_) );
  AD1V2C_8TH40 S2_2_11 ( .A(ab_2__11_), .B(n21), .CI(SUMB_1__12_), .CO(
        CARRYB_2__11_), .S(SUMB_2__11_) );
  AD1V2C_8TH40 S2_2_12 ( .A(ab_2__12_), .B(n20), .CI(SUMB_1__13_), .CO(
        CARRYB_2__12_), .S(SUMB_2__12_) );
  AD1V2C_8TH40 S2_2_13 ( .A(ab_2__13_), .B(n19), .CI(SUMB_1__14_), .CO(
        CARRYB_2__13_), .S(SUMB_2__13_) );
  AD1V2C_8TH40 S2_2_14 ( .A(ab_2__14_), .B(n18), .CI(SUMB_1__15_), .CO(
        CARRYB_2__14_), .S(SUMB_2__14_) );
  AD1V2C_8TH40 S2_2_15 ( .A(ab_2__15_), .B(n17), .CI(SUMB_1__16_), .CO(
        CARRYB_2__15_), .S(SUMB_2__15_) );
  AD1V2C_8TH40 S2_2_16 ( .A(ab_2__16_), .B(n16), .CI(SUMB_1__17_), .CO(
        CARRYB_2__16_), .S(SUMB_2__16_) );
  AD1V2C_8TH40 S2_2_17 ( .A(ab_2__17_), .B(n15), .CI(SUMB_1__18_), .CO(
        CARRYB_2__17_), .S(SUMB_2__17_) );
  AD1V2C_8TH40 S2_2_18 ( .A(ab_2__18_), .B(n14), .CI(SUMB_1__19_), .CO(
        CARRYB_2__18_), .S(SUMB_2__18_) );
  AD1V2C_8TH40 S2_2_19 ( .A(ab_2__19_), .B(n13), .CI(SUMB_1__20_), .CO(
        CARRYB_2__19_), .S(SUMB_2__19_) );
  AD1V2C_8TH40 S2_2_20 ( .A(ab_2__20_), .B(n12), .CI(SUMB_1__21_), .CO(
        CARRYB_2__20_), .S(SUMB_2__20_) );
  AD1V2C_8TH40 S2_2_21 ( .A(ab_2__21_), .B(n11), .CI(SUMB_1__22_), .CO(
        CARRYB_2__21_), .S(SUMB_2__21_) );
  AD1V2C_8TH40 S2_2_22 ( .A(ab_2__22_), .B(n10), .CI(SUMB_1__23_), .CO(
        CARRYB_2__22_), .S(SUMB_2__22_) );
  AD1V2C_8TH40 S2_2_23 ( .A(ab_2__23_), .B(n9), .CI(SUMB_1__24_), .CO(
        CARRYB_2__23_), .S(SUMB_2__23_) );
  AD1V2C_8TH40 S2_2_24 ( .A(ab_2__24_), .B(n8), .CI(SUMB_1__25_), .CO(
        CARRYB_2__24_), .S(SUMB_2__24_) );
  AD1V2C_8TH40 S2_2_25 ( .A(ab_2__25_), .B(n7), .CI(SUMB_1__26_), .CO(
        CARRYB_2__25_), .S(SUMB_2__25_) );
  AD1V2C_8TH40 S2_2_26 ( .A(ab_2__26_), .B(n6), .CI(SUMB_1__27_), .CO(
        CARRYB_2__26_), .S(SUMB_2__26_) );
  AD1V2C_8TH40 S2_2_27 ( .A(ab_2__27_), .B(n5), .CI(SUMB_1__28_), .CO(
        CARRYB_2__27_), .S(SUMB_2__27_) );
  AD1V2C_8TH40 S2_2_28 ( .A(ab_2__28_), .B(n4), .CI(SUMB_1__29_), .CO(
        CARRYB_2__28_), .S(SUMB_2__28_) );
  AD1V2C_8TH40 S2_2_29 ( .A(ab_2__29_), .B(n3), .CI(SUMB_1__30_), .CO(
        CARRYB_2__29_), .S(SUMB_2__29_) );
  AD1V2C_8TH40 S3_2_30 ( .A(ab_2__30_), .B(n2), .CI(ab_1__31_), .CO(
        CARRYB_2__30_), .S(SUMB_2__30_) );
  inst_execute_DW01_add_0 FS_1 ( .A({1'b0, A1_60_, A1_59_, A1_58_, A1_57_, 
        A1_56_, A1_55_, A1_54_, A1_53_, A1_52_, A1_51_, A1_50_, A1_49_, A1_48_, 
        A1_47_, A1_46_, A1_45_, A1_44_, A1_43_, A1_42_, A1_41_, A1_40_, A1_39_, 
        A1_38_, A1_37_, A1_36_, A1_35_, A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, 
        SUMB_31__0_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, 
        A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, 
        A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, 
        A1_3_, A1_2_, A1_1_, A1_0_}), .B({n33, n34, n57, n63, n56, n62, n55, 
        n61, n54, n60, n53, n59, n52, n58, n51, n50, n49, n48, n47, n46, n45, 
        n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[63:2]) );
  AND2V2_8TH40 U2 ( .A1(ab_1__30_), .A2(ab_0__31_), .Z(n2) );
  AND2V2_8TH40 U3 ( .A1(ab_1__29_), .A2(ab_0__30_), .Z(n3) );
  AND2V2_8TH40 U4 ( .A1(ab_1__28_), .A2(ab_0__29_), .Z(n4) );
  AND2V2_8TH40 U5 ( .A1(ab_1__27_), .A2(ab_0__28_), .Z(n5) );
  AND2V2_8TH40 U6 ( .A1(ab_1__26_), .A2(ab_0__27_), .Z(n6) );
  AND2V2_8TH40 U7 ( .A1(ab_1__25_), .A2(ab_0__26_), .Z(n7) );
  AND2V2_8TH40 U8 ( .A1(ab_1__24_), .A2(ab_0__25_), .Z(n8) );
  AND2V2_8TH40 U9 ( .A1(ab_1__23_), .A2(ab_0__24_), .Z(n9) );
  AND2V2_8TH40 U10 ( .A1(ab_1__22_), .A2(ab_0__23_), .Z(n10) );
  AND2V2_8TH40 U11 ( .A1(ab_1__21_), .A2(ab_0__22_), .Z(n11) );
  AND2V2_8TH40 U12 ( .A1(ab_1__20_), .A2(ab_0__21_), .Z(n12) );
  AND2V2_8TH40 U13 ( .A1(ab_1__19_), .A2(ab_0__20_), .Z(n13) );
  AND2V2_8TH40 U14 ( .A1(ab_1__18_), .A2(ab_0__19_), .Z(n14) );
  AND2V2_8TH40 U15 ( .A1(ab_1__17_), .A2(ab_0__18_), .Z(n15) );
  AND2V2_8TH40 U16 ( .A1(ab_1__16_), .A2(ab_0__17_), .Z(n16) );
  AND2V2_8TH40 U17 ( .A1(ab_1__15_), .A2(ab_0__16_), .Z(n17) );
  AND2V2_8TH40 U18 ( .A1(ab_1__14_), .A2(ab_0__15_), .Z(n18) );
  AND2V2_8TH40 U19 ( .A1(ab_1__13_), .A2(ab_0__14_), .Z(n19) );
  AND2V2_8TH40 U20 ( .A1(ab_1__12_), .A2(ab_0__13_), .Z(n20) );
  AND2V2_8TH40 U21 ( .A1(ab_1__11_), .A2(ab_0__12_), .Z(n21) );
  AND2V2_8TH40 U22 ( .A1(ab_1__10_), .A2(ab_0__11_), .Z(n22) );
  AND2V2_8TH40 U23 ( .A1(ab_1__9_), .A2(ab_0__10_), .Z(n23) );
  AND2V2_8TH40 U24 ( .A1(ab_1__8_), .A2(ab_0__9_), .Z(n24) );
  AND2V2_8TH40 U25 ( .A1(ab_1__7_), .A2(ab_0__8_), .Z(n25) );
  AND2V2_8TH40 U26 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(n26) );
  AND2V2_8TH40 U27 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(n27) );
  AND2V2_8TH40 U28 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(n28) );
  AND2V2_8TH40 U29 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(n29) );
  AND2V2_8TH40 U30 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(n30) );
  AND2V2_8TH40 U31 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(n31) );
  AND2V2_8TH40 U32 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(n32) );
  AND2V2_8TH40 U33 ( .A1(ab_31__31_), .A2(CARRYB_31__30_), .Z(n33) );
  AND2V2_8TH40 U34 ( .A1(SUMB_31__30_), .A2(CARRYB_31__29_), .Z(n34) );
  AND2V2_8TH40 U35 ( .A1(SUMB_31__1_), .A2(CARRYB_31__0_), .Z(n35) );
  AND2V2_8TH40 U36 ( .A1(SUMB_31__2_), .A2(CARRYB_31__1_), .Z(n36) );
  AND2V2_8TH40 U37 ( .A1(SUMB_31__3_), .A2(CARRYB_31__2_), .Z(n37) );
  AND2V2_8TH40 U38 ( .A1(SUMB_31__4_), .A2(CARRYB_31__3_), .Z(n38) );
  AND2V2_8TH40 U39 ( .A1(SUMB_31__5_), .A2(CARRYB_31__4_), .Z(n39) );
  AND2V2_8TH40 U40 ( .A1(SUMB_31__6_), .A2(CARRYB_31__5_), .Z(n40) );
  AND2V2_8TH40 U41 ( .A1(SUMB_31__7_), .A2(CARRYB_31__6_), .Z(n41) );
  AND2V2_8TH40 U42 ( .A1(SUMB_31__8_), .A2(CARRYB_31__7_), .Z(n42) );
  AND2V2_8TH40 U43 ( .A1(SUMB_31__9_), .A2(CARRYB_31__8_), .Z(n43) );
  AND2V2_8TH40 U44 ( .A1(SUMB_31__10_), .A2(CARRYB_31__9_), .Z(n44) );
  AND2V2_8TH40 U45 ( .A1(SUMB_31__11_), .A2(CARRYB_31__10_), .Z(n45) );
  AND2V2_8TH40 U46 ( .A1(SUMB_31__12_), .A2(CARRYB_31__11_), .Z(n46) );
  AND2V2_8TH40 U47 ( .A1(SUMB_31__13_), .A2(CARRYB_31__12_), .Z(n47) );
  AND2V2_8TH40 U48 ( .A1(SUMB_31__14_), .A2(CARRYB_31__13_), .Z(n48) );
  AND2V2_8TH40 U49 ( .A1(SUMB_31__15_), .A2(CARRYB_31__14_), .Z(n49) );
  AND2V2_8TH40 U50 ( .A1(SUMB_31__16_), .A2(CARRYB_31__15_), .Z(n50) );
  AND2V2_8TH40 U51 ( .A1(SUMB_31__17_), .A2(CARRYB_31__16_), .Z(n51) );
  AND2V2_8TH40 U52 ( .A1(SUMB_31__19_), .A2(CARRYB_31__18_), .Z(n52) );
  AND2V2_8TH40 U53 ( .A1(SUMB_31__21_), .A2(CARRYB_31__20_), .Z(n53) );
  AND2V2_8TH40 U54 ( .A1(SUMB_31__23_), .A2(CARRYB_31__22_), .Z(n54) );
  AND2V2_8TH40 U55 ( .A1(SUMB_31__25_), .A2(CARRYB_31__24_), .Z(n55) );
  AND2V2_8TH40 U56 ( .A1(SUMB_31__27_), .A2(CARRYB_31__26_), .Z(n56) );
  AND2V2_8TH40 U57 ( .A1(SUMB_31__29_), .A2(CARRYB_31__28_), .Z(n57) );
  AND2V2_8TH40 U58 ( .A1(SUMB_31__18_), .A2(CARRYB_31__17_), .Z(n58) );
  AND2V2_8TH40 U59 ( .A1(SUMB_31__20_), .A2(CARRYB_31__19_), .Z(n59) );
  AND2V2_8TH40 U60 ( .A1(SUMB_31__22_), .A2(CARRYB_31__21_), .Z(n60) );
  AND2V2_8TH40 U61 ( .A1(SUMB_31__24_), .A2(CARRYB_31__23_), .Z(n61) );
  AND2V2_8TH40 U62 ( .A1(SUMB_31__26_), .A2(CARRYB_31__25_), .Z(n62) );
  AND2V2_8TH40 U63 ( .A1(SUMB_31__28_), .A2(CARRYB_31__27_), .Z(n63) );
  INV2_8TH40 U64 ( .I(A[0]), .ZN(n64) );
  INV2_8TH40 U65 ( .I(A[3]), .ZN(n89) );
  INV2_8TH40 U66 ( .I(A[4]), .ZN(n90) );
  INV2_8TH40 U67 ( .I(A[5]), .ZN(n91) );
  INV2_8TH40 U68 ( .I(A[6]), .ZN(n92) );
  INV2_8TH40 U69 ( .I(A[7]), .ZN(n93) );
  INV2_8TH40 U70 ( .I(A[8]), .ZN(n94) );
  INV2_8TH40 U71 ( .I(A[10]), .ZN(n65) );
  INV2_8TH40 U72 ( .I(A[11]), .ZN(n66) );
  INV2_8TH40 U73 ( .I(A[2]), .ZN(n86) );
  INV2_8TH40 U74 ( .I(A[1]), .ZN(n75) );
  INV2_8TH40 U75 ( .I(A[12]), .ZN(n67) );
  INV2_8TH40 U76 ( .I(A[13]), .ZN(n68) );
  INV2_8TH40 U77 ( .I(A[14]), .ZN(n69) );
  INV2_8TH40 U78 ( .I(A[15]), .ZN(n70) );
  INV2_8TH40 U79 ( .I(A[16]), .ZN(n71) );
  INV2_8TH40 U80 ( .I(A[17]), .ZN(n72) );
  INV2_8TH40 U81 ( .I(A[18]), .ZN(n73) );
  INV2_8TH40 U82 ( .I(A[19]), .ZN(n74) );
  INV2_8TH40 U83 ( .I(A[20]), .ZN(n76) );
  INV2_8TH40 U84 ( .I(A[21]), .ZN(n77) );
  INV2_8TH40 U85 ( .I(A[22]), .ZN(n78) );
  INV2_8TH40 U86 ( .I(A[23]), .ZN(n79) );
  INV2_8TH40 U87 ( .I(A[24]), .ZN(n80) );
  INV2_8TH40 U88 ( .I(A[25]), .ZN(n81) );
  INV2_8TH40 U89 ( .I(A[26]), .ZN(n82) );
  INV2_8TH40 U90 ( .I(A[27]), .ZN(n83) );
  INV2_8TH40 U91 ( .I(A[28]), .ZN(n84) );
  INV2_8TH40 U92 ( .I(A[29]), .ZN(n85) );
  INV2_8TH40 U93 ( .I(A[30]), .ZN(n87) );
  INV2_8TH40 U94 ( .I(A[31]), .ZN(n88) );
  INV2_8TH40 U95 ( .I(B[0]), .ZN(n96) );
  INV2_8TH40 U96 ( .I(B[1]), .ZN(n107) );
  INV2_8TH40 U97 ( .I(B[2]), .ZN(n118) );
  INV2_8TH40 U98 ( .I(B[3]), .ZN(n121) );
  INV2_8TH40 U99 ( .I(B[4]), .ZN(n122) );
  INV2_8TH40 U100 ( .I(B[5]), .ZN(n123) );
  INV2_8TH40 U101 ( .I(B[6]), .ZN(n124) );
  INV2_8TH40 U102 ( .I(B[7]), .ZN(n125) );
  INV2_8TH40 U103 ( .I(B[8]), .ZN(n126) );
  INV2_8TH40 U104 ( .I(B[9]), .ZN(n127) );
  INV2_8TH40 U105 ( .I(B[10]), .ZN(n97) );
  INV2_8TH40 U106 ( .I(B[11]), .ZN(n98) );
  INV2_8TH40 U107 ( .I(B[12]), .ZN(n99) );
  INV2_8TH40 U108 ( .I(B[13]), .ZN(n100) );
  INV2_8TH40 U109 ( .I(B[14]), .ZN(n101) );
  INV2_8TH40 U110 ( .I(B[15]), .ZN(n102) );
  INV2_8TH40 U111 ( .I(B[16]), .ZN(n103) );
  INV2_8TH40 U112 ( .I(B[17]), .ZN(n104) );
  INV2_8TH40 U113 ( .I(B[18]), .ZN(n105) );
  INV2_8TH40 U114 ( .I(B[19]), .ZN(n106) );
  INV2_8TH40 U115 ( .I(B[20]), .ZN(n108) );
  INV2_8TH40 U116 ( .I(B[21]), .ZN(n109) );
  INV2_8TH40 U117 ( .I(B[24]), .ZN(n112) );
  INV2_8TH40 U118 ( .I(B[25]), .ZN(n113) );
  INV2_8TH40 U119 ( .I(B[23]), .ZN(n111) );
  INV2_8TH40 U120 ( .I(B[22]), .ZN(n110) );
  INV2_8TH40 U121 ( .I(B[26]), .ZN(n114) );
  INV2_8TH40 U122 ( .I(B[27]), .ZN(n115) );
  INV2_8TH40 U123 ( .I(B[28]), .ZN(n116) );
  INV2_8TH40 U124 ( .I(B[29]), .ZN(n117) );
  INV2_8TH40 U125 ( .I(B[30]), .ZN(n119) );
  INV2_8TH40 U126 ( .I(B[31]), .ZN(n120) );
  INV2_8TH40 U127 ( .I(A[9]), .ZN(n95) );
  XOR2V2_8TH40 U128 ( .A1(SUMB_31__1_), .A2(CARRYB_31__0_), .Z(A1_30_) );
  XOR2V2_8TH40 U129 ( .A1(SUMB_31__2_), .A2(CARRYB_31__1_), .Z(A1_31_) );
  XOR2V2_8TH40 U130 ( .A1(SUMB_31__3_), .A2(CARRYB_31__2_), .Z(A1_32_) );
  XOR2V2_8TH40 U131 ( .A1(SUMB_31__4_), .A2(CARRYB_31__3_), .Z(A1_33_) );
  XOR2V2_8TH40 U132 ( .A1(SUMB_31__5_), .A2(CARRYB_31__4_), .Z(A1_34_) );
  XOR2V2_8TH40 U133 ( .A1(SUMB_31__6_), .A2(CARRYB_31__5_), .Z(A1_35_) );
  XOR2V2_8TH40 U134 ( .A1(SUMB_31__7_), .A2(CARRYB_31__6_), .Z(A1_36_) );
  XOR2V2_8TH40 U135 ( .A1(SUMB_31__8_), .A2(CARRYB_31__7_), .Z(A1_37_) );
  XOR2V2_8TH40 U136 ( .A1(SUMB_31__9_), .A2(CARRYB_31__8_), .Z(A1_38_) );
  XOR2V2_8TH40 U137 ( .A1(SUMB_31__10_), .A2(CARRYB_31__9_), .Z(A1_39_) );
  XOR2V2_8TH40 U138 ( .A1(SUMB_31__11_), .A2(CARRYB_31__10_), .Z(A1_40_) );
  XOR2V2_8TH40 U139 ( .A1(SUMB_31__12_), .A2(CARRYB_31__11_), .Z(A1_41_) );
  XOR2V2_8TH40 U140 ( .A1(SUMB_31__13_), .A2(CARRYB_31__12_), .Z(A1_42_) );
  XOR2V2_8TH40 U141 ( .A1(SUMB_31__14_), .A2(CARRYB_31__13_), .Z(A1_43_) );
  XOR2V2_8TH40 U142 ( .A1(SUMB_31__15_), .A2(CARRYB_31__14_), .Z(A1_44_) );
  XOR2V2_8TH40 U143 ( .A1(SUMB_31__16_), .A2(CARRYB_31__15_), .Z(A1_45_) );
  XOR2V2_8TH40 U144 ( .A1(SUMB_31__17_), .A2(CARRYB_31__16_), .Z(A1_46_) );
  XOR2V2_8TH40 U145 ( .A1(SUMB_31__18_), .A2(CARRYB_31__17_), .Z(A1_47_) );
  XOR2V2_8TH40 U146 ( .A1(SUMB_31__19_), .A2(CARRYB_31__18_), .Z(A1_48_) );
  XOR2V2_8TH40 U147 ( .A1(SUMB_31__20_), .A2(CARRYB_31__19_), .Z(A1_49_) );
  XOR2V2_8TH40 U148 ( .A1(SUMB_31__21_), .A2(CARRYB_31__20_), .Z(A1_50_) );
  XOR2V2_8TH40 U149 ( .A1(SUMB_31__22_), .A2(CARRYB_31__21_), .Z(A1_51_) );
  XOR2V2_8TH40 U150 ( .A1(SUMB_31__23_), .A2(CARRYB_31__22_), .Z(A1_52_) );
  XOR2V2_8TH40 U151 ( .A1(SUMB_31__24_), .A2(CARRYB_31__23_), .Z(A1_53_) );
  XOR2V2_8TH40 U152 ( .A1(SUMB_31__25_), .A2(CARRYB_31__24_), .Z(A1_54_) );
  XOR2V2_8TH40 U153 ( .A1(SUMB_31__26_), .A2(CARRYB_31__25_), .Z(A1_55_) );
  XOR2V2_8TH40 U154 ( .A1(SUMB_31__27_), .A2(CARRYB_31__26_), .Z(A1_56_) );
  XOR2V2_8TH40 U155 ( .A1(SUMB_31__28_), .A2(CARRYB_31__27_), .Z(A1_57_) );
  XOR2V2_8TH40 U156 ( .A1(SUMB_31__29_), .A2(CARRYB_31__28_), .Z(A1_58_) );
  XOR2V2_8TH40 U157 ( .A1(SUMB_31__30_), .A2(CARRYB_31__29_), .Z(A1_59_) );
  XOR2V2_8TH40 U158 ( .A1(ab_31__31_), .A2(CARRYB_31__30_), .Z(A1_60_) );
  XOR2V2_8TH40 U159 ( .A1(ab_0__1_), .A2(ab_1__0_), .Z(PRODUCT[1]) );
  XOR2V2_8TH40 U160 ( .A1(ab_0__2_), .A2(ab_1__1_), .Z(SUMB_1__1_) );
  XOR2V2_8TH40 U161 ( .A1(ab_0__3_), .A2(ab_1__2_), .Z(SUMB_1__2_) );
  XOR2V2_8TH40 U162 ( .A1(ab_0__4_), .A2(ab_1__3_), .Z(SUMB_1__3_) );
  XOR2V2_8TH40 U163 ( .A1(ab_0__5_), .A2(ab_1__4_), .Z(SUMB_1__4_) );
  XOR2V2_8TH40 U164 ( .A1(ab_0__6_), .A2(ab_1__5_), .Z(SUMB_1__5_) );
  XOR2V2_8TH40 U165 ( .A1(ab_0__7_), .A2(ab_1__6_), .Z(SUMB_1__6_) );
  XOR2V2_8TH40 U166 ( .A1(ab_0__8_), .A2(ab_1__7_), .Z(SUMB_1__7_) );
  XOR2V2_8TH40 U167 ( .A1(ab_0__9_), .A2(ab_1__8_), .Z(SUMB_1__8_) );
  XOR2V2_8TH40 U168 ( .A1(ab_0__10_), .A2(ab_1__9_), .Z(SUMB_1__9_) );
  XOR2V2_8TH40 U169 ( .A1(ab_0__11_), .A2(ab_1__10_), .Z(SUMB_1__10_) );
  XOR2V2_8TH40 U170 ( .A1(ab_0__12_), .A2(ab_1__11_), .Z(SUMB_1__11_) );
  XOR2V2_8TH40 U171 ( .A1(ab_0__13_), .A2(ab_1__12_), .Z(SUMB_1__12_) );
  XOR2V2_8TH40 U172 ( .A1(ab_0__14_), .A2(ab_1__13_), .Z(SUMB_1__13_) );
  XOR2V2_8TH40 U173 ( .A1(ab_0__15_), .A2(ab_1__14_), .Z(SUMB_1__14_) );
  XOR2V2_8TH40 U174 ( .A1(ab_0__16_), .A2(ab_1__15_), .Z(SUMB_1__15_) );
  XOR2V2_8TH40 U175 ( .A1(ab_0__17_), .A2(ab_1__16_), .Z(SUMB_1__16_) );
  XOR2V2_8TH40 U176 ( .A1(ab_0__18_), .A2(ab_1__17_), .Z(SUMB_1__17_) );
  XOR2V2_8TH40 U177 ( .A1(ab_0__19_), .A2(ab_1__18_), .Z(SUMB_1__18_) );
  XOR2V2_8TH40 U178 ( .A1(ab_0__20_), .A2(ab_1__19_), .Z(SUMB_1__19_) );
  XOR2V2_8TH40 U179 ( .A1(ab_0__21_), .A2(ab_1__20_), .Z(SUMB_1__20_) );
  XOR2V2_8TH40 U180 ( .A1(ab_0__22_), .A2(ab_1__21_), .Z(SUMB_1__21_) );
  XOR2V2_8TH40 U181 ( .A1(ab_0__23_), .A2(ab_1__22_), .Z(SUMB_1__22_) );
  XOR2V2_8TH40 U182 ( .A1(ab_0__24_), .A2(ab_1__23_), .Z(SUMB_1__23_) );
  XOR2V2_8TH40 U183 ( .A1(ab_0__25_), .A2(ab_1__24_), .Z(SUMB_1__24_) );
  XOR2V2_8TH40 U184 ( .A1(ab_0__26_), .A2(ab_1__25_), .Z(SUMB_1__25_) );
  XOR2V2_8TH40 U185 ( .A1(ab_0__27_), .A2(ab_1__26_), .Z(SUMB_1__26_) );
  XOR2V2_8TH40 U186 ( .A1(ab_0__28_), .A2(ab_1__27_), .Z(SUMB_1__27_) );
  XOR2V2_8TH40 U187 ( .A1(ab_0__29_), .A2(ab_1__28_), .Z(SUMB_1__28_) );
  XOR2V2_8TH40 U188 ( .A1(ab_0__30_), .A2(ab_1__29_), .Z(SUMB_1__29_) );
  XOR2V2_8TH40 U189 ( .A1(ab_0__31_), .A2(ab_1__30_), .Z(SUMB_1__30_) );
  NOR2V0P5_8TH40 U191 ( .A1(n95), .A2(n127), .ZN(ab_9__9_) );
  NOR2V0P5_8TH40 U192 ( .A1(n95), .A2(n126), .ZN(ab_9__8_) );
  NOR2V0P5_8TH40 U193 ( .A1(n95), .A2(n125), .ZN(ab_9__7_) );
  NOR2V0P5_8TH40 U194 ( .A1(n95), .A2(n124), .ZN(ab_9__6_) );
  NOR2V0P5_8TH40 U195 ( .A1(n95), .A2(n123), .ZN(ab_9__5_) );
  NOR2V0P5_8TH40 U196 ( .A1(n95), .A2(n122), .ZN(ab_9__4_) );
  NOR2V0P5_8TH40 U197 ( .A1(n95), .A2(n121), .ZN(ab_9__3_) );
  NOR2V0P5_8TH40 U198 ( .A1(n95), .A2(n120), .ZN(ab_9__31_) );
  NOR2V0P5_8TH40 U199 ( .A1(n95), .A2(n119), .ZN(ab_9__30_) );
  NOR2V0P5_8TH40 U200 ( .A1(n95), .A2(n118), .ZN(ab_9__2_) );
  NOR2V0P5_8TH40 U201 ( .A1(n95), .A2(n117), .ZN(ab_9__29_) );
  NOR2V0P5_8TH40 U202 ( .A1(n95), .A2(n116), .ZN(ab_9__28_) );
  NOR2V0P5_8TH40 U203 ( .A1(n95), .A2(n115), .ZN(ab_9__27_) );
  NOR2V0P5_8TH40 U204 ( .A1(n95), .A2(n114), .ZN(ab_9__26_) );
  NOR2V0P5_8TH40 U205 ( .A1(n95), .A2(n113), .ZN(ab_9__25_) );
  NOR2V0P5_8TH40 U206 ( .A1(n95), .A2(n112), .ZN(ab_9__24_) );
  NOR2V0P5_8TH40 U207 ( .A1(n95), .A2(n111), .ZN(ab_9__23_) );
  NOR2V0P5_8TH40 U208 ( .A1(n95), .A2(n110), .ZN(ab_9__22_) );
  NOR2V0P5_8TH40 U209 ( .A1(n95), .A2(n109), .ZN(ab_9__21_) );
  NOR2V0P5_8TH40 U210 ( .A1(n95), .A2(n108), .ZN(ab_9__20_) );
  NOR2V0P5_8TH40 U211 ( .A1(n95), .A2(n107), .ZN(ab_9__1_) );
  NOR2V0P5_8TH40 U212 ( .A1(n95), .A2(n106), .ZN(ab_9__19_) );
  NOR2V0P5_8TH40 U213 ( .A1(n95), .A2(n105), .ZN(ab_9__18_) );
  NOR2V0P5_8TH40 U214 ( .A1(n95), .A2(n104), .ZN(ab_9__17_) );
  NOR2V0P5_8TH40 U215 ( .A1(n95), .A2(n103), .ZN(ab_9__16_) );
  NOR2V0P5_8TH40 U216 ( .A1(n95), .A2(n102), .ZN(ab_9__15_) );
  NOR2V0P5_8TH40 U217 ( .A1(n95), .A2(n101), .ZN(ab_9__14_) );
  NOR2V0P5_8TH40 U218 ( .A1(n95), .A2(n100), .ZN(ab_9__13_) );
  NOR2V0P5_8TH40 U219 ( .A1(n95), .A2(n99), .ZN(ab_9__12_) );
  NOR2V0P5_8TH40 U220 ( .A1(n95), .A2(n98), .ZN(ab_9__11_) );
  NOR2V0P5_8TH40 U221 ( .A1(n95), .A2(n97), .ZN(ab_9__10_) );
  NOR2V0P5_8TH40 U222 ( .A1(n95), .A2(n96), .ZN(ab_9__0_) );
  NOR2V0P5_8TH40 U223 ( .A1(n127), .A2(n94), .ZN(ab_8__9_) );
  NOR2V0P5_8TH40 U224 ( .A1(n126), .A2(n94), .ZN(ab_8__8_) );
  NOR2V0P5_8TH40 U225 ( .A1(n125), .A2(n94), .ZN(ab_8__7_) );
  NOR2V0P5_8TH40 U226 ( .A1(n124), .A2(n94), .ZN(ab_8__6_) );
  NOR2V0P5_8TH40 U227 ( .A1(n123), .A2(n94), .ZN(ab_8__5_) );
  NOR2V0P5_8TH40 U228 ( .A1(n122), .A2(n94), .ZN(ab_8__4_) );
  NOR2V0P5_8TH40 U229 ( .A1(n121), .A2(n94), .ZN(ab_8__3_) );
  NOR2V0P5_8TH40 U230 ( .A1(n120), .A2(n94), .ZN(ab_8__31_) );
  NOR2V0P5_8TH40 U231 ( .A1(n119), .A2(n94), .ZN(ab_8__30_) );
  NOR2V0P5_8TH40 U232 ( .A1(n118), .A2(n94), .ZN(ab_8__2_) );
  NOR2V0P5_8TH40 U233 ( .A1(n117), .A2(n94), .ZN(ab_8__29_) );
  NOR2V0P5_8TH40 U234 ( .A1(n116), .A2(n94), .ZN(ab_8__28_) );
  NOR2V0P5_8TH40 U235 ( .A1(n115), .A2(n94), .ZN(ab_8__27_) );
  NOR2V0P5_8TH40 U236 ( .A1(n114), .A2(n94), .ZN(ab_8__26_) );
  NOR2V0P5_8TH40 U237 ( .A1(n113), .A2(n94), .ZN(ab_8__25_) );
  NOR2V0P5_8TH40 U238 ( .A1(n112), .A2(n94), .ZN(ab_8__24_) );
  NOR2V0P5_8TH40 U239 ( .A1(n111), .A2(n94), .ZN(ab_8__23_) );
  NOR2V0P5_8TH40 U240 ( .A1(n110), .A2(n94), .ZN(ab_8__22_) );
  NOR2V0P5_8TH40 U241 ( .A1(n109), .A2(n94), .ZN(ab_8__21_) );
  NOR2V0P5_8TH40 U242 ( .A1(n108), .A2(n94), .ZN(ab_8__20_) );
  NOR2V0P5_8TH40 U243 ( .A1(n107), .A2(n94), .ZN(ab_8__1_) );
  NOR2V0P5_8TH40 U244 ( .A1(n106), .A2(n94), .ZN(ab_8__19_) );
  NOR2V0P5_8TH40 U245 ( .A1(n105), .A2(n94), .ZN(ab_8__18_) );
  NOR2V0P5_8TH40 U246 ( .A1(n104), .A2(n94), .ZN(ab_8__17_) );
  NOR2V0P5_8TH40 U247 ( .A1(n103), .A2(n94), .ZN(ab_8__16_) );
  NOR2V0P5_8TH40 U248 ( .A1(n102), .A2(n94), .ZN(ab_8__15_) );
  NOR2V0P5_8TH40 U249 ( .A1(n101), .A2(n94), .ZN(ab_8__14_) );
  NOR2V0P5_8TH40 U250 ( .A1(n100), .A2(n94), .ZN(ab_8__13_) );
  NOR2V0P5_8TH40 U251 ( .A1(n99), .A2(n94), .ZN(ab_8__12_) );
  NOR2V0P5_8TH40 U252 ( .A1(n98), .A2(n94), .ZN(ab_8__11_) );
  NOR2V0P5_8TH40 U253 ( .A1(n97), .A2(n94), .ZN(ab_8__10_) );
  NOR2V0P5_8TH40 U254 ( .A1(n96), .A2(n94), .ZN(ab_8__0_) );
  NOR2V0P5_8TH40 U255 ( .A1(n127), .A2(n93), .ZN(ab_7__9_) );
  NOR2V0P5_8TH40 U256 ( .A1(n126), .A2(n93), .ZN(ab_7__8_) );
  NOR2V0P5_8TH40 U257 ( .A1(n125), .A2(n93), .ZN(ab_7__7_) );
  NOR2V0P5_8TH40 U258 ( .A1(n124), .A2(n93), .ZN(ab_7__6_) );
  NOR2V0P5_8TH40 U259 ( .A1(n123), .A2(n93), .ZN(ab_7__5_) );
  NOR2V0P5_8TH40 U260 ( .A1(n122), .A2(n93), .ZN(ab_7__4_) );
  NOR2V0P5_8TH40 U261 ( .A1(n121), .A2(n93), .ZN(ab_7__3_) );
  NOR2V0P5_8TH40 U262 ( .A1(n120), .A2(n93), .ZN(ab_7__31_) );
  NOR2V0P5_8TH40 U263 ( .A1(n119), .A2(n93), .ZN(ab_7__30_) );
  NOR2V0P5_8TH40 U264 ( .A1(n118), .A2(n93), .ZN(ab_7__2_) );
  NOR2V0P5_8TH40 U265 ( .A1(n117), .A2(n93), .ZN(ab_7__29_) );
  NOR2V0P5_8TH40 U266 ( .A1(n116), .A2(n93), .ZN(ab_7__28_) );
  NOR2V0P5_8TH40 U267 ( .A1(n115), .A2(n93), .ZN(ab_7__27_) );
  NOR2V0P5_8TH40 U268 ( .A1(n114), .A2(n93), .ZN(ab_7__26_) );
  NOR2V0P5_8TH40 U269 ( .A1(n113), .A2(n93), .ZN(ab_7__25_) );
  NOR2V0P5_8TH40 U270 ( .A1(n112), .A2(n93), .ZN(ab_7__24_) );
  NOR2V0P5_8TH40 U271 ( .A1(n111), .A2(n93), .ZN(ab_7__23_) );
  NOR2V0P5_8TH40 U272 ( .A1(n110), .A2(n93), .ZN(ab_7__22_) );
  NOR2V0P5_8TH40 U273 ( .A1(n109), .A2(n93), .ZN(ab_7__21_) );
  NOR2V0P5_8TH40 U274 ( .A1(n108), .A2(n93), .ZN(ab_7__20_) );
  NOR2V0P5_8TH40 U275 ( .A1(n107), .A2(n93), .ZN(ab_7__1_) );
  NOR2V0P5_8TH40 U276 ( .A1(n106), .A2(n93), .ZN(ab_7__19_) );
  NOR2V0P5_8TH40 U277 ( .A1(n105), .A2(n93), .ZN(ab_7__18_) );
  NOR2V0P5_8TH40 U278 ( .A1(n104), .A2(n93), .ZN(ab_7__17_) );
  NOR2V0P5_8TH40 U279 ( .A1(n103), .A2(n93), .ZN(ab_7__16_) );
  NOR2V0P5_8TH40 U280 ( .A1(n102), .A2(n93), .ZN(ab_7__15_) );
  NOR2V0P5_8TH40 U281 ( .A1(n101), .A2(n93), .ZN(ab_7__14_) );
  NOR2V0P5_8TH40 U282 ( .A1(n100), .A2(n93), .ZN(ab_7__13_) );
  NOR2V0P5_8TH40 U283 ( .A1(n99), .A2(n93), .ZN(ab_7__12_) );
  NOR2V0P5_8TH40 U284 ( .A1(n98), .A2(n93), .ZN(ab_7__11_) );
  NOR2V0P5_8TH40 U285 ( .A1(n97), .A2(n93), .ZN(ab_7__10_) );
  NOR2V0P5_8TH40 U286 ( .A1(n96), .A2(n93), .ZN(ab_7__0_) );
  NOR2V0P5_8TH40 U287 ( .A1(n127), .A2(n92), .ZN(ab_6__9_) );
  NOR2V0P5_8TH40 U288 ( .A1(n126), .A2(n92), .ZN(ab_6__8_) );
  NOR2V0P5_8TH40 U289 ( .A1(n125), .A2(n92), .ZN(ab_6__7_) );
  NOR2V0P5_8TH40 U290 ( .A1(n124), .A2(n92), .ZN(ab_6__6_) );
  NOR2V0P5_8TH40 U291 ( .A1(n123), .A2(n92), .ZN(ab_6__5_) );
  NOR2V0P5_8TH40 U292 ( .A1(n122), .A2(n92), .ZN(ab_6__4_) );
  NOR2V0P5_8TH40 U293 ( .A1(n121), .A2(n92), .ZN(ab_6__3_) );
  NOR2V0P5_8TH40 U294 ( .A1(n120), .A2(n92), .ZN(ab_6__31_) );
  NOR2V0P5_8TH40 U295 ( .A1(n119), .A2(n92), .ZN(ab_6__30_) );
  NOR2V0P5_8TH40 U296 ( .A1(n118), .A2(n92), .ZN(ab_6__2_) );
  NOR2V0P5_8TH40 U297 ( .A1(n117), .A2(n92), .ZN(ab_6__29_) );
  NOR2V0P5_8TH40 U298 ( .A1(n116), .A2(n92), .ZN(ab_6__28_) );
  NOR2V0P5_8TH40 U299 ( .A1(n115), .A2(n92), .ZN(ab_6__27_) );
  NOR2V0P5_8TH40 U300 ( .A1(n114), .A2(n92), .ZN(ab_6__26_) );
  NOR2V0P5_8TH40 U301 ( .A1(n113), .A2(n92), .ZN(ab_6__25_) );
  NOR2V0P5_8TH40 U302 ( .A1(n112), .A2(n92), .ZN(ab_6__24_) );
  NOR2V0P5_8TH40 U303 ( .A1(n111), .A2(n92), .ZN(ab_6__23_) );
  NOR2V0P5_8TH40 U304 ( .A1(n110), .A2(n92), .ZN(ab_6__22_) );
  NOR2V0P5_8TH40 U305 ( .A1(n109), .A2(n92), .ZN(ab_6__21_) );
  NOR2V0P5_8TH40 U306 ( .A1(n108), .A2(n92), .ZN(ab_6__20_) );
  NOR2V0P5_8TH40 U307 ( .A1(n107), .A2(n92), .ZN(ab_6__1_) );
  NOR2V0P5_8TH40 U308 ( .A1(n106), .A2(n92), .ZN(ab_6__19_) );
  NOR2V0P5_8TH40 U309 ( .A1(n105), .A2(n92), .ZN(ab_6__18_) );
  NOR2V0P5_8TH40 U310 ( .A1(n104), .A2(n92), .ZN(ab_6__17_) );
  NOR2V0P5_8TH40 U311 ( .A1(n103), .A2(n92), .ZN(ab_6__16_) );
  NOR2V0P5_8TH40 U312 ( .A1(n102), .A2(n92), .ZN(ab_6__15_) );
  NOR2V0P5_8TH40 U313 ( .A1(n101), .A2(n92), .ZN(ab_6__14_) );
  NOR2V0P5_8TH40 U314 ( .A1(n100), .A2(n92), .ZN(ab_6__13_) );
  NOR2V0P5_8TH40 U315 ( .A1(n99), .A2(n92), .ZN(ab_6__12_) );
  NOR2V0P5_8TH40 U316 ( .A1(n98), .A2(n92), .ZN(ab_6__11_) );
  NOR2V0P5_8TH40 U317 ( .A1(n97), .A2(n92), .ZN(ab_6__10_) );
  NOR2V0P5_8TH40 U318 ( .A1(n96), .A2(n92), .ZN(ab_6__0_) );
  NOR2V0P5_8TH40 U319 ( .A1(n127), .A2(n91), .ZN(ab_5__9_) );
  NOR2V0P5_8TH40 U320 ( .A1(n126), .A2(n91), .ZN(ab_5__8_) );
  NOR2V0P5_8TH40 U321 ( .A1(n125), .A2(n91), .ZN(ab_5__7_) );
  NOR2V0P5_8TH40 U322 ( .A1(n124), .A2(n91), .ZN(ab_5__6_) );
  NOR2V0P5_8TH40 U323 ( .A1(n123), .A2(n91), .ZN(ab_5__5_) );
  NOR2V0P5_8TH40 U324 ( .A1(n122), .A2(n91), .ZN(ab_5__4_) );
  NOR2V0P5_8TH40 U325 ( .A1(n121), .A2(n91), .ZN(ab_5__3_) );
  NOR2V0P5_8TH40 U326 ( .A1(n120), .A2(n91), .ZN(ab_5__31_) );
  NOR2V0P5_8TH40 U327 ( .A1(n119), .A2(n91), .ZN(ab_5__30_) );
  NOR2V0P5_8TH40 U328 ( .A1(n118), .A2(n91), .ZN(ab_5__2_) );
  NOR2V0P5_8TH40 U329 ( .A1(n117), .A2(n91), .ZN(ab_5__29_) );
  NOR2V0P5_8TH40 U330 ( .A1(n116), .A2(n91), .ZN(ab_5__28_) );
  NOR2V0P5_8TH40 U331 ( .A1(n115), .A2(n91), .ZN(ab_5__27_) );
  NOR2V0P5_8TH40 U332 ( .A1(n114), .A2(n91), .ZN(ab_5__26_) );
  NOR2V0P5_8TH40 U333 ( .A1(n113), .A2(n91), .ZN(ab_5__25_) );
  NOR2V0P5_8TH40 U334 ( .A1(n112), .A2(n91), .ZN(ab_5__24_) );
  NOR2V0P5_8TH40 U335 ( .A1(n111), .A2(n91), .ZN(ab_5__23_) );
  NOR2V0P5_8TH40 U336 ( .A1(n110), .A2(n91), .ZN(ab_5__22_) );
  NOR2V0P5_8TH40 U337 ( .A1(n109), .A2(n91), .ZN(ab_5__21_) );
  NOR2V0P5_8TH40 U338 ( .A1(n108), .A2(n91), .ZN(ab_5__20_) );
  NOR2V0P5_8TH40 U339 ( .A1(n107), .A2(n91), .ZN(ab_5__1_) );
  NOR2V0P5_8TH40 U340 ( .A1(n106), .A2(n91), .ZN(ab_5__19_) );
  NOR2V0P5_8TH40 U341 ( .A1(n105), .A2(n91), .ZN(ab_5__18_) );
  NOR2V0P5_8TH40 U342 ( .A1(n104), .A2(n91), .ZN(ab_5__17_) );
  NOR2V0P5_8TH40 U343 ( .A1(n103), .A2(n91), .ZN(ab_5__16_) );
  NOR2V0P5_8TH40 U344 ( .A1(n102), .A2(n91), .ZN(ab_5__15_) );
  NOR2V0P5_8TH40 U345 ( .A1(n101), .A2(n91), .ZN(ab_5__14_) );
  NOR2V0P5_8TH40 U346 ( .A1(n100), .A2(n91), .ZN(ab_5__13_) );
  NOR2V0P5_8TH40 U347 ( .A1(n99), .A2(n91), .ZN(ab_5__12_) );
  NOR2V0P5_8TH40 U348 ( .A1(n98), .A2(n91), .ZN(ab_5__11_) );
  NOR2V0P5_8TH40 U349 ( .A1(n97), .A2(n91), .ZN(ab_5__10_) );
  NOR2V0P5_8TH40 U350 ( .A1(n96), .A2(n91), .ZN(ab_5__0_) );
  NOR2V0P5_8TH40 U351 ( .A1(n127), .A2(n90), .ZN(ab_4__9_) );
  NOR2V0P5_8TH40 U352 ( .A1(n126), .A2(n90), .ZN(ab_4__8_) );
  NOR2V0P5_8TH40 U353 ( .A1(n125), .A2(n90), .ZN(ab_4__7_) );
  NOR2V0P5_8TH40 U354 ( .A1(n124), .A2(n90), .ZN(ab_4__6_) );
  NOR2V0P5_8TH40 U355 ( .A1(n123), .A2(n90), .ZN(ab_4__5_) );
  NOR2V0P5_8TH40 U356 ( .A1(n122), .A2(n90), .ZN(ab_4__4_) );
  NOR2V0P5_8TH40 U357 ( .A1(n121), .A2(n90), .ZN(ab_4__3_) );
  NOR2V0P5_8TH40 U358 ( .A1(n120), .A2(n90), .ZN(ab_4__31_) );
  NOR2V0P5_8TH40 U359 ( .A1(n119), .A2(n90), .ZN(ab_4__30_) );
  NOR2V0P5_8TH40 U360 ( .A1(n118), .A2(n90), .ZN(ab_4__2_) );
  NOR2V0P5_8TH40 U361 ( .A1(n117), .A2(n90), .ZN(ab_4__29_) );
  NOR2V0P5_8TH40 U362 ( .A1(n116), .A2(n90), .ZN(ab_4__28_) );
  NOR2V0P5_8TH40 U363 ( .A1(n115), .A2(n90), .ZN(ab_4__27_) );
  NOR2V0P5_8TH40 U364 ( .A1(n114), .A2(n90), .ZN(ab_4__26_) );
  NOR2V0P5_8TH40 U365 ( .A1(n113), .A2(n90), .ZN(ab_4__25_) );
  NOR2V0P5_8TH40 U366 ( .A1(n112), .A2(n90), .ZN(ab_4__24_) );
  NOR2V0P5_8TH40 U367 ( .A1(n111), .A2(n90), .ZN(ab_4__23_) );
  NOR2V0P5_8TH40 U368 ( .A1(n110), .A2(n90), .ZN(ab_4__22_) );
  NOR2V0P5_8TH40 U369 ( .A1(n109), .A2(n90), .ZN(ab_4__21_) );
  NOR2V0P5_8TH40 U370 ( .A1(n108), .A2(n90), .ZN(ab_4__20_) );
  NOR2V0P5_8TH40 U371 ( .A1(n107), .A2(n90), .ZN(ab_4__1_) );
  NOR2V0P5_8TH40 U372 ( .A1(n106), .A2(n90), .ZN(ab_4__19_) );
  NOR2V0P5_8TH40 U373 ( .A1(n105), .A2(n90), .ZN(ab_4__18_) );
  NOR2V0P5_8TH40 U374 ( .A1(n104), .A2(n90), .ZN(ab_4__17_) );
  NOR2V0P5_8TH40 U375 ( .A1(n103), .A2(n90), .ZN(ab_4__16_) );
  NOR2V0P5_8TH40 U376 ( .A1(n102), .A2(n90), .ZN(ab_4__15_) );
  NOR2V0P5_8TH40 U377 ( .A1(n101), .A2(n90), .ZN(ab_4__14_) );
  NOR2V0P5_8TH40 U378 ( .A1(n100), .A2(n90), .ZN(ab_4__13_) );
  NOR2V0P5_8TH40 U379 ( .A1(n99), .A2(n90), .ZN(ab_4__12_) );
  NOR2V0P5_8TH40 U380 ( .A1(n98), .A2(n90), .ZN(ab_4__11_) );
  NOR2V0P5_8TH40 U381 ( .A1(n97), .A2(n90), .ZN(ab_4__10_) );
  NOR2V0P5_8TH40 U382 ( .A1(n96), .A2(n90), .ZN(ab_4__0_) );
  NOR2V0P5_8TH40 U383 ( .A1(n127), .A2(n89), .ZN(ab_3__9_) );
  NOR2V0P5_8TH40 U384 ( .A1(n126), .A2(n89), .ZN(ab_3__8_) );
  NOR2V0P5_8TH40 U385 ( .A1(n125), .A2(n89), .ZN(ab_3__7_) );
  NOR2V0P5_8TH40 U386 ( .A1(n124), .A2(n89), .ZN(ab_3__6_) );
  NOR2V0P5_8TH40 U387 ( .A1(n123), .A2(n89), .ZN(ab_3__5_) );
  NOR2V0P5_8TH40 U388 ( .A1(n122), .A2(n89), .ZN(ab_3__4_) );
  NOR2V0P5_8TH40 U389 ( .A1(n121), .A2(n89), .ZN(ab_3__3_) );
  NOR2V0P5_8TH40 U390 ( .A1(n120), .A2(n89), .ZN(ab_3__31_) );
  NOR2V0P5_8TH40 U391 ( .A1(n119), .A2(n89), .ZN(ab_3__30_) );
  NOR2V0P5_8TH40 U392 ( .A1(n118), .A2(n89), .ZN(ab_3__2_) );
  NOR2V0P5_8TH40 U393 ( .A1(n117), .A2(n89), .ZN(ab_3__29_) );
  NOR2V0P5_8TH40 U394 ( .A1(n116), .A2(n89), .ZN(ab_3__28_) );
  NOR2V0P5_8TH40 U395 ( .A1(n115), .A2(n89), .ZN(ab_3__27_) );
  NOR2V0P5_8TH40 U396 ( .A1(n114), .A2(n89), .ZN(ab_3__26_) );
  NOR2V0P5_8TH40 U397 ( .A1(n113), .A2(n89), .ZN(ab_3__25_) );
  NOR2V0P5_8TH40 U398 ( .A1(n112), .A2(n89), .ZN(ab_3__24_) );
  NOR2V0P5_8TH40 U399 ( .A1(n111), .A2(n89), .ZN(ab_3__23_) );
  NOR2V0P5_8TH40 U400 ( .A1(n110), .A2(n89), .ZN(ab_3__22_) );
  NOR2V0P5_8TH40 U401 ( .A1(n109), .A2(n89), .ZN(ab_3__21_) );
  NOR2V0P5_8TH40 U402 ( .A1(n108), .A2(n89), .ZN(ab_3__20_) );
  NOR2V0P5_8TH40 U403 ( .A1(n107), .A2(n89), .ZN(ab_3__1_) );
  NOR2V0P5_8TH40 U404 ( .A1(n106), .A2(n89), .ZN(ab_3__19_) );
  NOR2V0P5_8TH40 U405 ( .A1(n105), .A2(n89), .ZN(ab_3__18_) );
  NOR2V0P5_8TH40 U406 ( .A1(n104), .A2(n89), .ZN(ab_3__17_) );
  NOR2V0P5_8TH40 U407 ( .A1(n103), .A2(n89), .ZN(ab_3__16_) );
  NOR2V0P5_8TH40 U408 ( .A1(n102), .A2(n89), .ZN(ab_3__15_) );
  NOR2V0P5_8TH40 U409 ( .A1(n101), .A2(n89), .ZN(ab_3__14_) );
  NOR2V0P5_8TH40 U410 ( .A1(n100), .A2(n89), .ZN(ab_3__13_) );
  NOR2V0P5_8TH40 U411 ( .A1(n99), .A2(n89), .ZN(ab_3__12_) );
  NOR2V0P5_8TH40 U412 ( .A1(n98), .A2(n89), .ZN(ab_3__11_) );
  NOR2V0P5_8TH40 U413 ( .A1(n97), .A2(n89), .ZN(ab_3__10_) );
  NOR2V0P5_8TH40 U414 ( .A1(n96), .A2(n89), .ZN(ab_3__0_) );
  NOR2V0P5_8TH40 U415 ( .A1(n127), .A2(n88), .ZN(ab_31__9_) );
  NOR2V0P5_8TH40 U416 ( .A1(n126), .A2(n88), .ZN(ab_31__8_) );
  NOR2V0P5_8TH40 U417 ( .A1(n125), .A2(n88), .ZN(ab_31__7_) );
  NOR2V0P5_8TH40 U418 ( .A1(n124), .A2(n88), .ZN(ab_31__6_) );
  NOR2V0P5_8TH40 U419 ( .A1(n123), .A2(n88), .ZN(ab_31__5_) );
  NOR2V0P5_8TH40 U420 ( .A1(n122), .A2(n88), .ZN(ab_31__4_) );
  NOR2V0P5_8TH40 U421 ( .A1(n121), .A2(n88), .ZN(ab_31__3_) );
  NOR2V0P5_8TH40 U422 ( .A1(n120), .A2(n88), .ZN(ab_31__31_) );
  NOR2V0P5_8TH40 U423 ( .A1(n119), .A2(n88), .ZN(ab_31__30_) );
  NOR2V0P5_8TH40 U424 ( .A1(n118), .A2(n88), .ZN(ab_31__2_) );
  NOR2V0P5_8TH40 U425 ( .A1(n117), .A2(n88), .ZN(ab_31__29_) );
  NOR2V0P5_8TH40 U426 ( .A1(n116), .A2(n88), .ZN(ab_31__28_) );
  NOR2V0P5_8TH40 U427 ( .A1(n115), .A2(n88), .ZN(ab_31__27_) );
  NOR2V0P5_8TH40 U428 ( .A1(n114), .A2(n88), .ZN(ab_31__26_) );
  NOR2V0P5_8TH40 U429 ( .A1(n113), .A2(n88), .ZN(ab_31__25_) );
  NOR2V0P5_8TH40 U430 ( .A1(n112), .A2(n88), .ZN(ab_31__24_) );
  NOR2V0P5_8TH40 U431 ( .A1(n111), .A2(n88), .ZN(ab_31__23_) );
  NOR2V0P5_8TH40 U432 ( .A1(n110), .A2(n88), .ZN(ab_31__22_) );
  NOR2V0P5_8TH40 U433 ( .A1(n109), .A2(n88), .ZN(ab_31__21_) );
  NOR2V0P5_8TH40 U434 ( .A1(n108), .A2(n88), .ZN(ab_31__20_) );
  NOR2V0P5_8TH40 U435 ( .A1(n107), .A2(n88), .ZN(ab_31__1_) );
  NOR2V0P5_8TH40 U436 ( .A1(n106), .A2(n88), .ZN(ab_31__19_) );
  NOR2V0P5_8TH40 U437 ( .A1(n105), .A2(n88), .ZN(ab_31__18_) );
  NOR2V0P5_8TH40 U438 ( .A1(n104), .A2(n88), .ZN(ab_31__17_) );
  NOR2V0P5_8TH40 U439 ( .A1(n103), .A2(n88), .ZN(ab_31__16_) );
  NOR2V0P5_8TH40 U440 ( .A1(n102), .A2(n88), .ZN(ab_31__15_) );
  NOR2V0P5_8TH40 U441 ( .A1(n101), .A2(n88), .ZN(ab_31__14_) );
  NOR2V0P5_8TH40 U442 ( .A1(n100), .A2(n88), .ZN(ab_31__13_) );
  NOR2V0P5_8TH40 U443 ( .A1(n99), .A2(n88), .ZN(ab_31__12_) );
  NOR2V0P5_8TH40 U444 ( .A1(n98), .A2(n88), .ZN(ab_31__11_) );
  NOR2V0P5_8TH40 U445 ( .A1(n97), .A2(n88), .ZN(ab_31__10_) );
  NOR2V0P5_8TH40 U446 ( .A1(n96), .A2(n88), .ZN(ab_31__0_) );
  NOR2V0P5_8TH40 U447 ( .A1(n127), .A2(n87), .ZN(ab_30__9_) );
  NOR2V0P5_8TH40 U448 ( .A1(n126), .A2(n87), .ZN(ab_30__8_) );
  NOR2V0P5_8TH40 U449 ( .A1(n125), .A2(n87), .ZN(ab_30__7_) );
  NOR2V0P5_8TH40 U450 ( .A1(n124), .A2(n87), .ZN(ab_30__6_) );
  NOR2V0P5_8TH40 U451 ( .A1(n123), .A2(n87), .ZN(ab_30__5_) );
  NOR2V0P5_8TH40 U452 ( .A1(n122), .A2(n87), .ZN(ab_30__4_) );
  NOR2V0P5_8TH40 U453 ( .A1(n121), .A2(n87), .ZN(ab_30__3_) );
  NOR2V0P5_8TH40 U454 ( .A1(n120), .A2(n87), .ZN(ab_30__31_) );
  NOR2V0P5_8TH40 U455 ( .A1(n119), .A2(n87), .ZN(ab_30__30_) );
  NOR2V0P5_8TH40 U456 ( .A1(n118), .A2(n87), .ZN(ab_30__2_) );
  NOR2V0P5_8TH40 U457 ( .A1(n117), .A2(n87), .ZN(ab_30__29_) );
  NOR2V0P5_8TH40 U458 ( .A1(n116), .A2(n87), .ZN(ab_30__28_) );
  NOR2V0P5_8TH40 U459 ( .A1(n115), .A2(n87), .ZN(ab_30__27_) );
  NOR2V0P5_8TH40 U460 ( .A1(n114), .A2(n87), .ZN(ab_30__26_) );
  NOR2V0P5_8TH40 U461 ( .A1(n113), .A2(n87), .ZN(ab_30__25_) );
  NOR2V0P5_8TH40 U462 ( .A1(n112), .A2(n87), .ZN(ab_30__24_) );
  NOR2V0P5_8TH40 U463 ( .A1(n111), .A2(n87), .ZN(ab_30__23_) );
  NOR2V0P5_8TH40 U464 ( .A1(n110), .A2(n87), .ZN(ab_30__22_) );
  NOR2V0P5_8TH40 U465 ( .A1(n109), .A2(n87), .ZN(ab_30__21_) );
  NOR2V0P5_8TH40 U466 ( .A1(n108), .A2(n87), .ZN(ab_30__20_) );
  NOR2V0P5_8TH40 U467 ( .A1(n107), .A2(n87), .ZN(ab_30__1_) );
  NOR2V0P5_8TH40 U468 ( .A1(n106), .A2(n87), .ZN(ab_30__19_) );
  NOR2V0P5_8TH40 U469 ( .A1(n105), .A2(n87), .ZN(ab_30__18_) );
  NOR2V0P5_8TH40 U470 ( .A1(n104), .A2(n87), .ZN(ab_30__17_) );
  NOR2V0P5_8TH40 U471 ( .A1(n103), .A2(n87), .ZN(ab_30__16_) );
  NOR2V0P5_8TH40 U472 ( .A1(n102), .A2(n87), .ZN(ab_30__15_) );
  NOR2V0P5_8TH40 U473 ( .A1(n101), .A2(n87), .ZN(ab_30__14_) );
  NOR2V0P5_8TH40 U474 ( .A1(n100), .A2(n87), .ZN(ab_30__13_) );
  NOR2V0P5_8TH40 U475 ( .A1(n99), .A2(n87), .ZN(ab_30__12_) );
  NOR2V0P5_8TH40 U476 ( .A1(n98), .A2(n87), .ZN(ab_30__11_) );
  NOR2V0P5_8TH40 U477 ( .A1(n97), .A2(n87), .ZN(ab_30__10_) );
  NOR2V0P5_8TH40 U478 ( .A1(n96), .A2(n87), .ZN(ab_30__0_) );
  NOR2V0P5_8TH40 U479 ( .A1(n127), .A2(n86), .ZN(ab_2__9_) );
  NOR2V0P5_8TH40 U480 ( .A1(n126), .A2(n86), .ZN(ab_2__8_) );
  NOR2V0P5_8TH40 U481 ( .A1(n125), .A2(n86), .ZN(ab_2__7_) );
  NOR2V0P5_8TH40 U482 ( .A1(n124), .A2(n86), .ZN(ab_2__6_) );
  NOR2V0P5_8TH40 U483 ( .A1(n123), .A2(n86), .ZN(ab_2__5_) );
  NOR2V0P5_8TH40 U484 ( .A1(n122), .A2(n86), .ZN(ab_2__4_) );
  NOR2V0P5_8TH40 U485 ( .A1(n121), .A2(n86), .ZN(ab_2__3_) );
  NOR2V0P5_8TH40 U486 ( .A1(n120), .A2(n86), .ZN(ab_2__31_) );
  NOR2V0P5_8TH40 U487 ( .A1(n119), .A2(n86), .ZN(ab_2__30_) );
  NOR2V0P5_8TH40 U488 ( .A1(n118), .A2(n86), .ZN(ab_2__2_) );
  NOR2V0P5_8TH40 U489 ( .A1(n117), .A2(n86), .ZN(ab_2__29_) );
  NOR2V0P5_8TH40 U490 ( .A1(n116), .A2(n86), .ZN(ab_2__28_) );
  NOR2V0P5_8TH40 U491 ( .A1(n115), .A2(n86), .ZN(ab_2__27_) );
  NOR2V0P5_8TH40 U492 ( .A1(n114), .A2(n86), .ZN(ab_2__26_) );
  NOR2V0P5_8TH40 U493 ( .A1(n113), .A2(n86), .ZN(ab_2__25_) );
  NOR2V0P5_8TH40 U494 ( .A1(n112), .A2(n86), .ZN(ab_2__24_) );
  NOR2V0P5_8TH40 U495 ( .A1(n111), .A2(n86), .ZN(ab_2__23_) );
  NOR2V0P5_8TH40 U496 ( .A1(n110), .A2(n86), .ZN(ab_2__22_) );
  NOR2V0P5_8TH40 U497 ( .A1(n109), .A2(n86), .ZN(ab_2__21_) );
  NOR2V0P5_8TH40 U498 ( .A1(n108), .A2(n86), .ZN(ab_2__20_) );
  NOR2V0P5_8TH40 U499 ( .A1(n107), .A2(n86), .ZN(ab_2__1_) );
  NOR2V0P5_8TH40 U500 ( .A1(n106), .A2(n86), .ZN(ab_2__19_) );
  NOR2V0P5_8TH40 U501 ( .A1(n105), .A2(n86), .ZN(ab_2__18_) );
  NOR2V0P5_8TH40 U502 ( .A1(n104), .A2(n86), .ZN(ab_2__17_) );
  NOR2V0P5_8TH40 U503 ( .A1(n103), .A2(n86), .ZN(ab_2__16_) );
  NOR2V0P5_8TH40 U504 ( .A1(n102), .A2(n86), .ZN(ab_2__15_) );
  NOR2V0P5_8TH40 U505 ( .A1(n101), .A2(n86), .ZN(ab_2__14_) );
  NOR2V0P5_8TH40 U506 ( .A1(n100), .A2(n86), .ZN(ab_2__13_) );
  NOR2V0P5_8TH40 U507 ( .A1(n99), .A2(n86), .ZN(ab_2__12_) );
  NOR2V0P5_8TH40 U508 ( .A1(n98), .A2(n86), .ZN(ab_2__11_) );
  NOR2V0P5_8TH40 U509 ( .A1(n97), .A2(n86), .ZN(ab_2__10_) );
  NOR2V0P5_8TH40 U510 ( .A1(n96), .A2(n86), .ZN(ab_2__0_) );
  NOR2V0P5_8TH40 U511 ( .A1(n127), .A2(n85), .ZN(ab_29__9_) );
  NOR2V0P5_8TH40 U512 ( .A1(n126), .A2(n85), .ZN(ab_29__8_) );
  NOR2V0P5_8TH40 U513 ( .A1(n125), .A2(n85), .ZN(ab_29__7_) );
  NOR2V0P5_8TH40 U514 ( .A1(n124), .A2(n85), .ZN(ab_29__6_) );
  NOR2V0P5_8TH40 U515 ( .A1(n123), .A2(n85), .ZN(ab_29__5_) );
  NOR2V0P5_8TH40 U516 ( .A1(n122), .A2(n85), .ZN(ab_29__4_) );
  NOR2V0P5_8TH40 U517 ( .A1(n121), .A2(n85), .ZN(ab_29__3_) );
  NOR2V0P5_8TH40 U518 ( .A1(n120), .A2(n85), .ZN(ab_29__31_) );
  NOR2V0P5_8TH40 U519 ( .A1(n119), .A2(n85), .ZN(ab_29__30_) );
  NOR2V0P5_8TH40 U520 ( .A1(n118), .A2(n85), .ZN(ab_29__2_) );
  NOR2V0P5_8TH40 U521 ( .A1(n117), .A2(n85), .ZN(ab_29__29_) );
  NOR2V0P5_8TH40 U522 ( .A1(n116), .A2(n85), .ZN(ab_29__28_) );
  NOR2V0P5_8TH40 U523 ( .A1(n115), .A2(n85), .ZN(ab_29__27_) );
  NOR2V0P5_8TH40 U524 ( .A1(n114), .A2(n85), .ZN(ab_29__26_) );
  NOR2V0P5_8TH40 U525 ( .A1(n113), .A2(n85), .ZN(ab_29__25_) );
  NOR2V0P5_8TH40 U526 ( .A1(n112), .A2(n85), .ZN(ab_29__24_) );
  NOR2V0P5_8TH40 U527 ( .A1(n111), .A2(n85), .ZN(ab_29__23_) );
  NOR2V0P5_8TH40 U528 ( .A1(n110), .A2(n85), .ZN(ab_29__22_) );
  NOR2V0P5_8TH40 U529 ( .A1(n109), .A2(n85), .ZN(ab_29__21_) );
  NOR2V0P5_8TH40 U530 ( .A1(n108), .A2(n85), .ZN(ab_29__20_) );
  NOR2V0P5_8TH40 U531 ( .A1(n107), .A2(n85), .ZN(ab_29__1_) );
  NOR2V0P5_8TH40 U532 ( .A1(n106), .A2(n85), .ZN(ab_29__19_) );
  NOR2V0P5_8TH40 U533 ( .A1(n105), .A2(n85), .ZN(ab_29__18_) );
  NOR2V0P5_8TH40 U534 ( .A1(n104), .A2(n85), .ZN(ab_29__17_) );
  NOR2V0P5_8TH40 U535 ( .A1(n103), .A2(n85), .ZN(ab_29__16_) );
  NOR2V0P5_8TH40 U536 ( .A1(n102), .A2(n85), .ZN(ab_29__15_) );
  NOR2V0P5_8TH40 U537 ( .A1(n101), .A2(n85), .ZN(ab_29__14_) );
  NOR2V0P5_8TH40 U538 ( .A1(n100), .A2(n85), .ZN(ab_29__13_) );
  NOR2V0P5_8TH40 U539 ( .A1(n99), .A2(n85), .ZN(ab_29__12_) );
  NOR2V0P5_8TH40 U540 ( .A1(n98), .A2(n85), .ZN(ab_29__11_) );
  NOR2V0P5_8TH40 U541 ( .A1(n97), .A2(n85), .ZN(ab_29__10_) );
  NOR2V0P5_8TH40 U542 ( .A1(n96), .A2(n85), .ZN(ab_29__0_) );
  NOR2V0P5_8TH40 U543 ( .A1(n127), .A2(n84), .ZN(ab_28__9_) );
  NOR2V0P5_8TH40 U544 ( .A1(n126), .A2(n84), .ZN(ab_28__8_) );
  NOR2V0P5_8TH40 U545 ( .A1(n125), .A2(n84), .ZN(ab_28__7_) );
  NOR2V0P5_8TH40 U546 ( .A1(n124), .A2(n84), .ZN(ab_28__6_) );
  NOR2V0P5_8TH40 U547 ( .A1(n123), .A2(n84), .ZN(ab_28__5_) );
  NOR2V0P5_8TH40 U548 ( .A1(n122), .A2(n84), .ZN(ab_28__4_) );
  NOR2V0P5_8TH40 U549 ( .A1(n121), .A2(n84), .ZN(ab_28__3_) );
  NOR2V0P5_8TH40 U550 ( .A1(n120), .A2(n84), .ZN(ab_28__31_) );
  NOR2V0P5_8TH40 U551 ( .A1(n119), .A2(n84), .ZN(ab_28__30_) );
  NOR2V0P5_8TH40 U552 ( .A1(n118), .A2(n84), .ZN(ab_28__2_) );
  NOR2V0P5_8TH40 U553 ( .A1(n117), .A2(n84), .ZN(ab_28__29_) );
  NOR2V0P5_8TH40 U554 ( .A1(n116), .A2(n84), .ZN(ab_28__28_) );
  NOR2V0P5_8TH40 U555 ( .A1(n115), .A2(n84), .ZN(ab_28__27_) );
  NOR2V0P5_8TH40 U556 ( .A1(n114), .A2(n84), .ZN(ab_28__26_) );
  NOR2V0P5_8TH40 U557 ( .A1(n113), .A2(n84), .ZN(ab_28__25_) );
  NOR2V0P5_8TH40 U558 ( .A1(n112), .A2(n84), .ZN(ab_28__24_) );
  NOR2V0P5_8TH40 U559 ( .A1(n111), .A2(n84), .ZN(ab_28__23_) );
  NOR2V0P5_8TH40 U560 ( .A1(n110), .A2(n84), .ZN(ab_28__22_) );
  NOR2V0P5_8TH40 U561 ( .A1(n109), .A2(n84), .ZN(ab_28__21_) );
  NOR2V0P5_8TH40 U562 ( .A1(n108), .A2(n84), .ZN(ab_28__20_) );
  NOR2V0P5_8TH40 U563 ( .A1(n107), .A2(n84), .ZN(ab_28__1_) );
  NOR2V0P5_8TH40 U564 ( .A1(n106), .A2(n84), .ZN(ab_28__19_) );
  NOR2V0P5_8TH40 U565 ( .A1(n105), .A2(n84), .ZN(ab_28__18_) );
  NOR2V0P5_8TH40 U566 ( .A1(n104), .A2(n84), .ZN(ab_28__17_) );
  NOR2V0P5_8TH40 U567 ( .A1(n103), .A2(n84), .ZN(ab_28__16_) );
  NOR2V0P5_8TH40 U568 ( .A1(n102), .A2(n84), .ZN(ab_28__15_) );
  NOR2V0P5_8TH40 U569 ( .A1(n101), .A2(n84), .ZN(ab_28__14_) );
  NOR2V0P5_8TH40 U570 ( .A1(n100), .A2(n84), .ZN(ab_28__13_) );
  NOR2V0P5_8TH40 U571 ( .A1(n99), .A2(n84), .ZN(ab_28__12_) );
  NOR2V0P5_8TH40 U572 ( .A1(n98), .A2(n84), .ZN(ab_28__11_) );
  NOR2V0P5_8TH40 U573 ( .A1(n97), .A2(n84), .ZN(ab_28__10_) );
  NOR2V0P5_8TH40 U574 ( .A1(n96), .A2(n84), .ZN(ab_28__0_) );
  NOR2V0P5_8TH40 U575 ( .A1(n127), .A2(n83), .ZN(ab_27__9_) );
  NOR2V0P5_8TH40 U576 ( .A1(n126), .A2(n83), .ZN(ab_27__8_) );
  NOR2V0P5_8TH40 U577 ( .A1(n125), .A2(n83), .ZN(ab_27__7_) );
  NOR2V0P5_8TH40 U578 ( .A1(n124), .A2(n83), .ZN(ab_27__6_) );
  NOR2V0P5_8TH40 U579 ( .A1(n123), .A2(n83), .ZN(ab_27__5_) );
  NOR2V0P5_8TH40 U580 ( .A1(n122), .A2(n83), .ZN(ab_27__4_) );
  NOR2V0P5_8TH40 U581 ( .A1(n121), .A2(n83), .ZN(ab_27__3_) );
  NOR2V0P5_8TH40 U582 ( .A1(n120), .A2(n83), .ZN(ab_27__31_) );
  NOR2V0P5_8TH40 U583 ( .A1(n119), .A2(n83), .ZN(ab_27__30_) );
  NOR2V0P5_8TH40 U584 ( .A1(n118), .A2(n83), .ZN(ab_27__2_) );
  NOR2V0P5_8TH40 U585 ( .A1(n117), .A2(n83), .ZN(ab_27__29_) );
  NOR2V0P5_8TH40 U586 ( .A1(n116), .A2(n83), .ZN(ab_27__28_) );
  NOR2V0P5_8TH40 U587 ( .A1(n115), .A2(n83), .ZN(ab_27__27_) );
  NOR2V0P5_8TH40 U588 ( .A1(n114), .A2(n83), .ZN(ab_27__26_) );
  NOR2V0P5_8TH40 U589 ( .A1(n113), .A2(n83), .ZN(ab_27__25_) );
  NOR2V0P5_8TH40 U590 ( .A1(n112), .A2(n83), .ZN(ab_27__24_) );
  NOR2V0P5_8TH40 U591 ( .A1(n111), .A2(n83), .ZN(ab_27__23_) );
  NOR2V0P5_8TH40 U592 ( .A1(n110), .A2(n83), .ZN(ab_27__22_) );
  NOR2V0P5_8TH40 U593 ( .A1(n109), .A2(n83), .ZN(ab_27__21_) );
  NOR2V0P5_8TH40 U594 ( .A1(n108), .A2(n83), .ZN(ab_27__20_) );
  NOR2V0P5_8TH40 U595 ( .A1(n107), .A2(n83), .ZN(ab_27__1_) );
  NOR2V0P5_8TH40 U596 ( .A1(n106), .A2(n83), .ZN(ab_27__19_) );
  NOR2V0P5_8TH40 U597 ( .A1(n105), .A2(n83), .ZN(ab_27__18_) );
  NOR2V0P5_8TH40 U598 ( .A1(n104), .A2(n83), .ZN(ab_27__17_) );
  NOR2V0P5_8TH40 U599 ( .A1(n103), .A2(n83), .ZN(ab_27__16_) );
  NOR2V0P5_8TH40 U600 ( .A1(n102), .A2(n83), .ZN(ab_27__15_) );
  NOR2V0P5_8TH40 U601 ( .A1(n101), .A2(n83), .ZN(ab_27__14_) );
  NOR2V0P5_8TH40 U602 ( .A1(n100), .A2(n83), .ZN(ab_27__13_) );
  NOR2V0P5_8TH40 U603 ( .A1(n99), .A2(n83), .ZN(ab_27__12_) );
  NOR2V0P5_8TH40 U604 ( .A1(n98), .A2(n83), .ZN(ab_27__11_) );
  NOR2V0P5_8TH40 U605 ( .A1(n97), .A2(n83), .ZN(ab_27__10_) );
  NOR2V0P5_8TH40 U606 ( .A1(n96), .A2(n83), .ZN(ab_27__0_) );
  NOR2V0P5_8TH40 U607 ( .A1(n127), .A2(n82), .ZN(ab_26__9_) );
  NOR2V0P5_8TH40 U608 ( .A1(n126), .A2(n82), .ZN(ab_26__8_) );
  NOR2V0P5_8TH40 U609 ( .A1(n125), .A2(n82), .ZN(ab_26__7_) );
  NOR2V0P5_8TH40 U610 ( .A1(n124), .A2(n82), .ZN(ab_26__6_) );
  NOR2V0P5_8TH40 U611 ( .A1(n123), .A2(n82), .ZN(ab_26__5_) );
  NOR2V0P5_8TH40 U612 ( .A1(n122), .A2(n82), .ZN(ab_26__4_) );
  NOR2V0P5_8TH40 U613 ( .A1(n121), .A2(n82), .ZN(ab_26__3_) );
  NOR2V0P5_8TH40 U614 ( .A1(n120), .A2(n82), .ZN(ab_26__31_) );
  NOR2V0P5_8TH40 U615 ( .A1(n119), .A2(n82), .ZN(ab_26__30_) );
  NOR2V0P5_8TH40 U616 ( .A1(n118), .A2(n82), .ZN(ab_26__2_) );
  NOR2V0P5_8TH40 U617 ( .A1(n117), .A2(n82), .ZN(ab_26__29_) );
  NOR2V0P5_8TH40 U618 ( .A1(n116), .A2(n82), .ZN(ab_26__28_) );
  NOR2V0P5_8TH40 U619 ( .A1(n115), .A2(n82), .ZN(ab_26__27_) );
  NOR2V0P5_8TH40 U620 ( .A1(n114), .A2(n82), .ZN(ab_26__26_) );
  NOR2V0P5_8TH40 U621 ( .A1(n113), .A2(n82), .ZN(ab_26__25_) );
  NOR2V0P5_8TH40 U622 ( .A1(n112), .A2(n82), .ZN(ab_26__24_) );
  NOR2V0P5_8TH40 U623 ( .A1(n111), .A2(n82), .ZN(ab_26__23_) );
  NOR2V0P5_8TH40 U624 ( .A1(n110), .A2(n82), .ZN(ab_26__22_) );
  NOR2V0P5_8TH40 U625 ( .A1(n109), .A2(n82), .ZN(ab_26__21_) );
  NOR2V0P5_8TH40 U626 ( .A1(n108), .A2(n82), .ZN(ab_26__20_) );
  NOR2V0P5_8TH40 U627 ( .A1(n107), .A2(n82), .ZN(ab_26__1_) );
  NOR2V0P5_8TH40 U628 ( .A1(n106), .A2(n82), .ZN(ab_26__19_) );
  NOR2V0P5_8TH40 U629 ( .A1(n105), .A2(n82), .ZN(ab_26__18_) );
  NOR2V0P5_8TH40 U630 ( .A1(n104), .A2(n82), .ZN(ab_26__17_) );
  NOR2V0P5_8TH40 U631 ( .A1(n103), .A2(n82), .ZN(ab_26__16_) );
  NOR2V0P5_8TH40 U632 ( .A1(n102), .A2(n82), .ZN(ab_26__15_) );
  NOR2V0P5_8TH40 U633 ( .A1(n101), .A2(n82), .ZN(ab_26__14_) );
  NOR2V0P5_8TH40 U634 ( .A1(n100), .A2(n82), .ZN(ab_26__13_) );
  NOR2V0P5_8TH40 U635 ( .A1(n99), .A2(n82), .ZN(ab_26__12_) );
  NOR2V0P5_8TH40 U636 ( .A1(n98), .A2(n82), .ZN(ab_26__11_) );
  NOR2V0P5_8TH40 U637 ( .A1(n97), .A2(n82), .ZN(ab_26__10_) );
  NOR2V0P5_8TH40 U638 ( .A1(n96), .A2(n82), .ZN(ab_26__0_) );
  NOR2V0P5_8TH40 U639 ( .A1(n127), .A2(n81), .ZN(ab_25__9_) );
  NOR2V0P5_8TH40 U640 ( .A1(n126), .A2(n81), .ZN(ab_25__8_) );
  NOR2V0P5_8TH40 U641 ( .A1(n125), .A2(n81), .ZN(ab_25__7_) );
  NOR2V0P5_8TH40 U642 ( .A1(n124), .A2(n81), .ZN(ab_25__6_) );
  NOR2V0P5_8TH40 U643 ( .A1(n123), .A2(n81), .ZN(ab_25__5_) );
  NOR2V0P5_8TH40 U644 ( .A1(n122), .A2(n81), .ZN(ab_25__4_) );
  NOR2V0P5_8TH40 U645 ( .A1(n121), .A2(n81), .ZN(ab_25__3_) );
  NOR2V0P5_8TH40 U646 ( .A1(n120), .A2(n81), .ZN(ab_25__31_) );
  NOR2V0P5_8TH40 U647 ( .A1(n119), .A2(n81), .ZN(ab_25__30_) );
  NOR2V0P5_8TH40 U648 ( .A1(n118), .A2(n81), .ZN(ab_25__2_) );
  NOR2V0P5_8TH40 U649 ( .A1(n117), .A2(n81), .ZN(ab_25__29_) );
  NOR2V0P5_8TH40 U650 ( .A1(n116), .A2(n81), .ZN(ab_25__28_) );
  NOR2V0P5_8TH40 U651 ( .A1(n115), .A2(n81), .ZN(ab_25__27_) );
  NOR2V0P5_8TH40 U652 ( .A1(n114), .A2(n81), .ZN(ab_25__26_) );
  NOR2V0P5_8TH40 U653 ( .A1(n113), .A2(n81), .ZN(ab_25__25_) );
  NOR2V0P5_8TH40 U654 ( .A1(n112), .A2(n81), .ZN(ab_25__24_) );
  NOR2V0P5_8TH40 U655 ( .A1(n111), .A2(n81), .ZN(ab_25__23_) );
  NOR2V0P5_8TH40 U656 ( .A1(n110), .A2(n81), .ZN(ab_25__22_) );
  NOR2V0P5_8TH40 U657 ( .A1(n109), .A2(n81), .ZN(ab_25__21_) );
  NOR2V0P5_8TH40 U658 ( .A1(n108), .A2(n81), .ZN(ab_25__20_) );
  NOR2V0P5_8TH40 U659 ( .A1(n107), .A2(n81), .ZN(ab_25__1_) );
  NOR2V0P5_8TH40 U660 ( .A1(n106), .A2(n81), .ZN(ab_25__19_) );
  NOR2V0P5_8TH40 U661 ( .A1(n105), .A2(n81), .ZN(ab_25__18_) );
  NOR2V0P5_8TH40 U662 ( .A1(n104), .A2(n81), .ZN(ab_25__17_) );
  NOR2V0P5_8TH40 U663 ( .A1(n103), .A2(n81), .ZN(ab_25__16_) );
  NOR2V0P5_8TH40 U664 ( .A1(n102), .A2(n81), .ZN(ab_25__15_) );
  NOR2V0P5_8TH40 U665 ( .A1(n101), .A2(n81), .ZN(ab_25__14_) );
  NOR2V0P5_8TH40 U666 ( .A1(n100), .A2(n81), .ZN(ab_25__13_) );
  NOR2V0P5_8TH40 U667 ( .A1(n99), .A2(n81), .ZN(ab_25__12_) );
  NOR2V0P5_8TH40 U668 ( .A1(n98), .A2(n81), .ZN(ab_25__11_) );
  NOR2V0P5_8TH40 U669 ( .A1(n97), .A2(n81), .ZN(ab_25__10_) );
  NOR2V0P5_8TH40 U670 ( .A1(n96), .A2(n81), .ZN(ab_25__0_) );
  NOR2V0P5_8TH40 U671 ( .A1(n127), .A2(n80), .ZN(ab_24__9_) );
  NOR2V0P5_8TH40 U672 ( .A1(n126), .A2(n80), .ZN(ab_24__8_) );
  NOR2V0P5_8TH40 U673 ( .A1(n125), .A2(n80), .ZN(ab_24__7_) );
  NOR2V0P5_8TH40 U674 ( .A1(n124), .A2(n80), .ZN(ab_24__6_) );
  NOR2V0P5_8TH40 U675 ( .A1(n123), .A2(n80), .ZN(ab_24__5_) );
  NOR2V0P5_8TH40 U676 ( .A1(n122), .A2(n80), .ZN(ab_24__4_) );
  NOR2V0P5_8TH40 U677 ( .A1(n121), .A2(n80), .ZN(ab_24__3_) );
  NOR2V0P5_8TH40 U678 ( .A1(n120), .A2(n80), .ZN(ab_24__31_) );
  NOR2V0P5_8TH40 U679 ( .A1(n119), .A2(n80), .ZN(ab_24__30_) );
  NOR2V0P5_8TH40 U680 ( .A1(n118), .A2(n80), .ZN(ab_24__2_) );
  NOR2V0P5_8TH40 U681 ( .A1(n117), .A2(n80), .ZN(ab_24__29_) );
  NOR2V0P5_8TH40 U682 ( .A1(n116), .A2(n80), .ZN(ab_24__28_) );
  NOR2V0P5_8TH40 U683 ( .A1(n115), .A2(n80), .ZN(ab_24__27_) );
  NOR2V0P5_8TH40 U684 ( .A1(n114), .A2(n80), .ZN(ab_24__26_) );
  NOR2V0P5_8TH40 U685 ( .A1(n113), .A2(n80), .ZN(ab_24__25_) );
  NOR2V0P5_8TH40 U686 ( .A1(n112), .A2(n80), .ZN(ab_24__24_) );
  NOR2V0P5_8TH40 U687 ( .A1(n111), .A2(n80), .ZN(ab_24__23_) );
  NOR2V0P5_8TH40 U688 ( .A1(n110), .A2(n80), .ZN(ab_24__22_) );
  NOR2V0P5_8TH40 U689 ( .A1(n109), .A2(n80), .ZN(ab_24__21_) );
  NOR2V0P5_8TH40 U690 ( .A1(n108), .A2(n80), .ZN(ab_24__20_) );
  NOR2V0P5_8TH40 U691 ( .A1(n107), .A2(n80), .ZN(ab_24__1_) );
  NOR2V0P5_8TH40 U692 ( .A1(n106), .A2(n80), .ZN(ab_24__19_) );
  NOR2V0P5_8TH40 U693 ( .A1(n105), .A2(n80), .ZN(ab_24__18_) );
  NOR2V0P5_8TH40 U694 ( .A1(n104), .A2(n80), .ZN(ab_24__17_) );
  NOR2V0P5_8TH40 U695 ( .A1(n103), .A2(n80), .ZN(ab_24__16_) );
  NOR2V0P5_8TH40 U696 ( .A1(n102), .A2(n80), .ZN(ab_24__15_) );
  NOR2V0P5_8TH40 U697 ( .A1(n101), .A2(n80), .ZN(ab_24__14_) );
  NOR2V0P5_8TH40 U698 ( .A1(n100), .A2(n80), .ZN(ab_24__13_) );
  NOR2V0P5_8TH40 U699 ( .A1(n99), .A2(n80), .ZN(ab_24__12_) );
  NOR2V0P5_8TH40 U700 ( .A1(n98), .A2(n80), .ZN(ab_24__11_) );
  NOR2V0P5_8TH40 U701 ( .A1(n97), .A2(n80), .ZN(ab_24__10_) );
  NOR2V0P5_8TH40 U702 ( .A1(n96), .A2(n80), .ZN(ab_24__0_) );
  NOR2V0P5_8TH40 U703 ( .A1(n127), .A2(n79), .ZN(ab_23__9_) );
  NOR2V0P5_8TH40 U704 ( .A1(n126), .A2(n79), .ZN(ab_23__8_) );
  NOR2V0P5_8TH40 U705 ( .A1(n125), .A2(n79), .ZN(ab_23__7_) );
  NOR2V0P5_8TH40 U706 ( .A1(n124), .A2(n79), .ZN(ab_23__6_) );
  NOR2V0P5_8TH40 U707 ( .A1(n123), .A2(n79), .ZN(ab_23__5_) );
  NOR2V0P5_8TH40 U708 ( .A1(n122), .A2(n79), .ZN(ab_23__4_) );
  NOR2V0P5_8TH40 U709 ( .A1(n121), .A2(n79), .ZN(ab_23__3_) );
  NOR2V0P5_8TH40 U710 ( .A1(n120), .A2(n79), .ZN(ab_23__31_) );
  NOR2V0P5_8TH40 U711 ( .A1(n119), .A2(n79), .ZN(ab_23__30_) );
  NOR2V0P5_8TH40 U712 ( .A1(n118), .A2(n79), .ZN(ab_23__2_) );
  NOR2V0P5_8TH40 U713 ( .A1(n117), .A2(n79), .ZN(ab_23__29_) );
  NOR2V0P5_8TH40 U714 ( .A1(n116), .A2(n79), .ZN(ab_23__28_) );
  NOR2V0P5_8TH40 U715 ( .A1(n115), .A2(n79), .ZN(ab_23__27_) );
  NOR2V0P5_8TH40 U716 ( .A1(n114), .A2(n79), .ZN(ab_23__26_) );
  NOR2V0P5_8TH40 U717 ( .A1(n113), .A2(n79), .ZN(ab_23__25_) );
  NOR2V0P5_8TH40 U718 ( .A1(n112), .A2(n79), .ZN(ab_23__24_) );
  NOR2V0P5_8TH40 U719 ( .A1(n111), .A2(n79), .ZN(ab_23__23_) );
  NOR2V0P5_8TH40 U720 ( .A1(n110), .A2(n79), .ZN(ab_23__22_) );
  NOR2V0P5_8TH40 U721 ( .A1(n109), .A2(n79), .ZN(ab_23__21_) );
  NOR2V0P5_8TH40 U722 ( .A1(n108), .A2(n79), .ZN(ab_23__20_) );
  NOR2V0P5_8TH40 U723 ( .A1(n107), .A2(n79), .ZN(ab_23__1_) );
  NOR2V0P5_8TH40 U724 ( .A1(n106), .A2(n79), .ZN(ab_23__19_) );
  NOR2V0P5_8TH40 U725 ( .A1(n105), .A2(n79), .ZN(ab_23__18_) );
  NOR2V0P5_8TH40 U726 ( .A1(n104), .A2(n79), .ZN(ab_23__17_) );
  NOR2V0P5_8TH40 U727 ( .A1(n103), .A2(n79), .ZN(ab_23__16_) );
  NOR2V0P5_8TH40 U728 ( .A1(n102), .A2(n79), .ZN(ab_23__15_) );
  NOR2V0P5_8TH40 U729 ( .A1(n101), .A2(n79), .ZN(ab_23__14_) );
  NOR2V0P5_8TH40 U730 ( .A1(n100), .A2(n79), .ZN(ab_23__13_) );
  NOR2V0P5_8TH40 U731 ( .A1(n99), .A2(n79), .ZN(ab_23__12_) );
  NOR2V0P5_8TH40 U732 ( .A1(n98), .A2(n79), .ZN(ab_23__11_) );
  NOR2V0P5_8TH40 U733 ( .A1(n97), .A2(n79), .ZN(ab_23__10_) );
  NOR2V0P5_8TH40 U734 ( .A1(n96), .A2(n79), .ZN(ab_23__0_) );
  NOR2V0P5_8TH40 U735 ( .A1(n127), .A2(n78), .ZN(ab_22__9_) );
  NOR2V0P5_8TH40 U736 ( .A1(n126), .A2(n78), .ZN(ab_22__8_) );
  NOR2V0P5_8TH40 U737 ( .A1(n125), .A2(n78), .ZN(ab_22__7_) );
  NOR2V0P5_8TH40 U738 ( .A1(n124), .A2(n78), .ZN(ab_22__6_) );
  NOR2V0P5_8TH40 U739 ( .A1(n123), .A2(n78), .ZN(ab_22__5_) );
  NOR2V0P5_8TH40 U740 ( .A1(n122), .A2(n78), .ZN(ab_22__4_) );
  NOR2V0P5_8TH40 U741 ( .A1(n121), .A2(n78), .ZN(ab_22__3_) );
  NOR2V0P5_8TH40 U742 ( .A1(n120), .A2(n78), .ZN(ab_22__31_) );
  NOR2V0P5_8TH40 U743 ( .A1(n119), .A2(n78), .ZN(ab_22__30_) );
  NOR2V0P5_8TH40 U744 ( .A1(n118), .A2(n78), .ZN(ab_22__2_) );
  NOR2V0P5_8TH40 U745 ( .A1(n117), .A2(n78), .ZN(ab_22__29_) );
  NOR2V0P5_8TH40 U746 ( .A1(n116), .A2(n78), .ZN(ab_22__28_) );
  NOR2V0P5_8TH40 U747 ( .A1(n115), .A2(n78), .ZN(ab_22__27_) );
  NOR2V0P5_8TH40 U748 ( .A1(n114), .A2(n78), .ZN(ab_22__26_) );
  NOR2V0P5_8TH40 U749 ( .A1(n113), .A2(n78), .ZN(ab_22__25_) );
  NOR2V0P5_8TH40 U750 ( .A1(n112), .A2(n78), .ZN(ab_22__24_) );
  NOR2V0P5_8TH40 U751 ( .A1(n111), .A2(n78), .ZN(ab_22__23_) );
  NOR2V0P5_8TH40 U752 ( .A1(n110), .A2(n78), .ZN(ab_22__22_) );
  NOR2V0P5_8TH40 U753 ( .A1(n109), .A2(n78), .ZN(ab_22__21_) );
  NOR2V0P5_8TH40 U754 ( .A1(n108), .A2(n78), .ZN(ab_22__20_) );
  NOR2V0P5_8TH40 U755 ( .A1(n107), .A2(n78), .ZN(ab_22__1_) );
  NOR2V0P5_8TH40 U756 ( .A1(n106), .A2(n78), .ZN(ab_22__19_) );
  NOR2V0P5_8TH40 U757 ( .A1(n105), .A2(n78), .ZN(ab_22__18_) );
  NOR2V0P5_8TH40 U758 ( .A1(n104), .A2(n78), .ZN(ab_22__17_) );
  NOR2V0P5_8TH40 U759 ( .A1(n103), .A2(n78), .ZN(ab_22__16_) );
  NOR2V0P5_8TH40 U760 ( .A1(n102), .A2(n78), .ZN(ab_22__15_) );
  NOR2V0P5_8TH40 U761 ( .A1(n101), .A2(n78), .ZN(ab_22__14_) );
  NOR2V0P5_8TH40 U762 ( .A1(n100), .A2(n78), .ZN(ab_22__13_) );
  NOR2V0P5_8TH40 U763 ( .A1(n99), .A2(n78), .ZN(ab_22__12_) );
  NOR2V0P5_8TH40 U764 ( .A1(n98), .A2(n78), .ZN(ab_22__11_) );
  NOR2V0P5_8TH40 U765 ( .A1(n97), .A2(n78), .ZN(ab_22__10_) );
  NOR2V0P5_8TH40 U766 ( .A1(n96), .A2(n78), .ZN(ab_22__0_) );
  NOR2V0P5_8TH40 U767 ( .A1(n127), .A2(n77), .ZN(ab_21__9_) );
  NOR2V0P5_8TH40 U768 ( .A1(n126), .A2(n77), .ZN(ab_21__8_) );
  NOR2V0P5_8TH40 U769 ( .A1(n125), .A2(n77), .ZN(ab_21__7_) );
  NOR2V0P5_8TH40 U770 ( .A1(n124), .A2(n77), .ZN(ab_21__6_) );
  NOR2V0P5_8TH40 U771 ( .A1(n123), .A2(n77), .ZN(ab_21__5_) );
  NOR2V0P5_8TH40 U772 ( .A1(n122), .A2(n77), .ZN(ab_21__4_) );
  NOR2V0P5_8TH40 U773 ( .A1(n121), .A2(n77), .ZN(ab_21__3_) );
  NOR2V0P5_8TH40 U774 ( .A1(n120), .A2(n77), .ZN(ab_21__31_) );
  NOR2V0P5_8TH40 U775 ( .A1(n119), .A2(n77), .ZN(ab_21__30_) );
  NOR2V0P5_8TH40 U776 ( .A1(n118), .A2(n77), .ZN(ab_21__2_) );
  NOR2V0P5_8TH40 U777 ( .A1(n117), .A2(n77), .ZN(ab_21__29_) );
  NOR2V0P5_8TH40 U778 ( .A1(n116), .A2(n77), .ZN(ab_21__28_) );
  NOR2V0P5_8TH40 U779 ( .A1(n115), .A2(n77), .ZN(ab_21__27_) );
  NOR2V0P5_8TH40 U780 ( .A1(n114), .A2(n77), .ZN(ab_21__26_) );
  NOR2V0P5_8TH40 U781 ( .A1(n113), .A2(n77), .ZN(ab_21__25_) );
  NOR2V0P5_8TH40 U782 ( .A1(n112), .A2(n77), .ZN(ab_21__24_) );
  NOR2V0P5_8TH40 U783 ( .A1(n111), .A2(n77), .ZN(ab_21__23_) );
  NOR2V0P5_8TH40 U784 ( .A1(n110), .A2(n77), .ZN(ab_21__22_) );
  NOR2V0P5_8TH40 U785 ( .A1(n109), .A2(n77), .ZN(ab_21__21_) );
  NOR2V0P5_8TH40 U786 ( .A1(n108), .A2(n77), .ZN(ab_21__20_) );
  NOR2V0P5_8TH40 U787 ( .A1(n107), .A2(n77), .ZN(ab_21__1_) );
  NOR2V0P5_8TH40 U788 ( .A1(n106), .A2(n77), .ZN(ab_21__19_) );
  NOR2V0P5_8TH40 U789 ( .A1(n105), .A2(n77), .ZN(ab_21__18_) );
  NOR2V0P5_8TH40 U790 ( .A1(n104), .A2(n77), .ZN(ab_21__17_) );
  NOR2V0P5_8TH40 U791 ( .A1(n103), .A2(n77), .ZN(ab_21__16_) );
  NOR2V0P5_8TH40 U792 ( .A1(n102), .A2(n77), .ZN(ab_21__15_) );
  NOR2V0P5_8TH40 U793 ( .A1(n101), .A2(n77), .ZN(ab_21__14_) );
  NOR2V0P5_8TH40 U794 ( .A1(n100), .A2(n77), .ZN(ab_21__13_) );
  NOR2V0P5_8TH40 U795 ( .A1(n99), .A2(n77), .ZN(ab_21__12_) );
  NOR2V0P5_8TH40 U796 ( .A1(n98), .A2(n77), .ZN(ab_21__11_) );
  NOR2V0P5_8TH40 U797 ( .A1(n97), .A2(n77), .ZN(ab_21__10_) );
  NOR2V0P5_8TH40 U798 ( .A1(n96), .A2(n77), .ZN(ab_21__0_) );
  NOR2V0P5_8TH40 U799 ( .A1(n127), .A2(n76), .ZN(ab_20__9_) );
  NOR2V0P5_8TH40 U800 ( .A1(n126), .A2(n76), .ZN(ab_20__8_) );
  NOR2V0P5_8TH40 U801 ( .A1(n125), .A2(n76), .ZN(ab_20__7_) );
  NOR2V0P5_8TH40 U802 ( .A1(n124), .A2(n76), .ZN(ab_20__6_) );
  NOR2V0P5_8TH40 U803 ( .A1(n123), .A2(n76), .ZN(ab_20__5_) );
  NOR2V0P5_8TH40 U804 ( .A1(n122), .A2(n76), .ZN(ab_20__4_) );
  NOR2V0P5_8TH40 U805 ( .A1(n121), .A2(n76), .ZN(ab_20__3_) );
  NOR2V0P5_8TH40 U806 ( .A1(n120), .A2(n76), .ZN(ab_20__31_) );
  NOR2V0P5_8TH40 U807 ( .A1(n119), .A2(n76), .ZN(ab_20__30_) );
  NOR2V0P5_8TH40 U808 ( .A1(n118), .A2(n76), .ZN(ab_20__2_) );
  NOR2V0P5_8TH40 U809 ( .A1(n117), .A2(n76), .ZN(ab_20__29_) );
  NOR2V0P5_8TH40 U810 ( .A1(n116), .A2(n76), .ZN(ab_20__28_) );
  NOR2V0P5_8TH40 U811 ( .A1(n115), .A2(n76), .ZN(ab_20__27_) );
  NOR2V0P5_8TH40 U812 ( .A1(n114), .A2(n76), .ZN(ab_20__26_) );
  NOR2V0P5_8TH40 U813 ( .A1(n113), .A2(n76), .ZN(ab_20__25_) );
  NOR2V0P5_8TH40 U814 ( .A1(n112), .A2(n76), .ZN(ab_20__24_) );
  NOR2V0P5_8TH40 U815 ( .A1(n111), .A2(n76), .ZN(ab_20__23_) );
  NOR2V0P5_8TH40 U816 ( .A1(n110), .A2(n76), .ZN(ab_20__22_) );
  NOR2V0P5_8TH40 U817 ( .A1(n109), .A2(n76), .ZN(ab_20__21_) );
  NOR2V0P5_8TH40 U818 ( .A1(n108), .A2(n76), .ZN(ab_20__20_) );
  NOR2V0P5_8TH40 U819 ( .A1(n107), .A2(n76), .ZN(ab_20__1_) );
  NOR2V0P5_8TH40 U820 ( .A1(n106), .A2(n76), .ZN(ab_20__19_) );
  NOR2V0P5_8TH40 U821 ( .A1(n105), .A2(n76), .ZN(ab_20__18_) );
  NOR2V0P5_8TH40 U822 ( .A1(n104), .A2(n76), .ZN(ab_20__17_) );
  NOR2V0P5_8TH40 U823 ( .A1(n103), .A2(n76), .ZN(ab_20__16_) );
  NOR2V0P5_8TH40 U824 ( .A1(n102), .A2(n76), .ZN(ab_20__15_) );
  NOR2V0P5_8TH40 U825 ( .A1(n101), .A2(n76), .ZN(ab_20__14_) );
  NOR2V0P5_8TH40 U826 ( .A1(n100), .A2(n76), .ZN(ab_20__13_) );
  NOR2V0P5_8TH40 U827 ( .A1(n99), .A2(n76), .ZN(ab_20__12_) );
  NOR2V0P5_8TH40 U828 ( .A1(n98), .A2(n76), .ZN(ab_20__11_) );
  NOR2V0P5_8TH40 U829 ( .A1(n97), .A2(n76), .ZN(ab_20__10_) );
  NOR2V0P5_8TH40 U830 ( .A1(n96), .A2(n76), .ZN(ab_20__0_) );
  NOR2V0P5_8TH40 U831 ( .A1(n127), .A2(n75), .ZN(ab_1__9_) );
  NOR2V0P5_8TH40 U832 ( .A1(n126), .A2(n75), .ZN(ab_1__8_) );
  NOR2V0P5_8TH40 U833 ( .A1(n125), .A2(n75), .ZN(ab_1__7_) );
  NOR2V0P5_8TH40 U834 ( .A1(n124), .A2(n75), .ZN(ab_1__6_) );
  NOR2V0P5_8TH40 U835 ( .A1(n123), .A2(n75), .ZN(ab_1__5_) );
  NOR2V0P5_8TH40 U836 ( .A1(n122), .A2(n75), .ZN(ab_1__4_) );
  NOR2V0P5_8TH40 U837 ( .A1(n121), .A2(n75), .ZN(ab_1__3_) );
  NOR2V0P5_8TH40 U838 ( .A1(n120), .A2(n75), .ZN(ab_1__31_) );
  NOR2V0P5_8TH40 U839 ( .A1(n119), .A2(n75), .ZN(ab_1__30_) );
  NOR2V0P5_8TH40 U840 ( .A1(n118), .A2(n75), .ZN(ab_1__2_) );
  NOR2V0P5_8TH40 U841 ( .A1(n117), .A2(n75), .ZN(ab_1__29_) );
  NOR2V0P5_8TH40 U842 ( .A1(n116), .A2(n75), .ZN(ab_1__28_) );
  NOR2V0P5_8TH40 U843 ( .A1(n115), .A2(n75), .ZN(ab_1__27_) );
  NOR2V0P5_8TH40 U844 ( .A1(n114), .A2(n75), .ZN(ab_1__26_) );
  NOR2V0P5_8TH40 U845 ( .A1(n113), .A2(n75), .ZN(ab_1__25_) );
  NOR2V0P5_8TH40 U846 ( .A1(n112), .A2(n75), .ZN(ab_1__24_) );
  NOR2V0P5_8TH40 U847 ( .A1(n111), .A2(n75), .ZN(ab_1__23_) );
  NOR2V0P5_8TH40 U848 ( .A1(n110), .A2(n75), .ZN(ab_1__22_) );
  NOR2V0P5_8TH40 U849 ( .A1(n109), .A2(n75), .ZN(ab_1__21_) );
  NOR2V0P5_8TH40 U850 ( .A1(n108), .A2(n75), .ZN(ab_1__20_) );
  NOR2V0P5_8TH40 U851 ( .A1(n107), .A2(n75), .ZN(ab_1__1_) );
  NOR2V0P5_8TH40 U852 ( .A1(n106), .A2(n75), .ZN(ab_1__19_) );
  NOR2V0P5_8TH40 U853 ( .A1(n105), .A2(n75), .ZN(ab_1__18_) );
  NOR2V0P5_8TH40 U854 ( .A1(n104), .A2(n75), .ZN(ab_1__17_) );
  NOR2V0P5_8TH40 U855 ( .A1(n103), .A2(n75), .ZN(ab_1__16_) );
  NOR2V0P5_8TH40 U856 ( .A1(n102), .A2(n75), .ZN(ab_1__15_) );
  NOR2V0P5_8TH40 U857 ( .A1(n101), .A2(n75), .ZN(ab_1__14_) );
  NOR2V0P5_8TH40 U858 ( .A1(n100), .A2(n75), .ZN(ab_1__13_) );
  NOR2V0P5_8TH40 U859 ( .A1(n99), .A2(n75), .ZN(ab_1__12_) );
  NOR2V0P5_8TH40 U860 ( .A1(n98), .A2(n75), .ZN(ab_1__11_) );
  NOR2V0P5_8TH40 U861 ( .A1(n97), .A2(n75), .ZN(ab_1__10_) );
  NOR2V0P5_8TH40 U862 ( .A1(n96), .A2(n75), .ZN(ab_1__0_) );
  NOR2V0P5_8TH40 U863 ( .A1(n127), .A2(n74), .ZN(ab_19__9_) );
  NOR2V0P5_8TH40 U864 ( .A1(n126), .A2(n74), .ZN(ab_19__8_) );
  NOR2V0P5_8TH40 U865 ( .A1(n125), .A2(n74), .ZN(ab_19__7_) );
  NOR2V0P5_8TH40 U866 ( .A1(n124), .A2(n74), .ZN(ab_19__6_) );
  NOR2V0P5_8TH40 U867 ( .A1(n123), .A2(n74), .ZN(ab_19__5_) );
  NOR2V0P5_8TH40 U868 ( .A1(n122), .A2(n74), .ZN(ab_19__4_) );
  NOR2V0P5_8TH40 U869 ( .A1(n121), .A2(n74), .ZN(ab_19__3_) );
  NOR2V0P5_8TH40 U870 ( .A1(n120), .A2(n74), .ZN(ab_19__31_) );
  NOR2V0P5_8TH40 U871 ( .A1(n119), .A2(n74), .ZN(ab_19__30_) );
  NOR2V0P5_8TH40 U872 ( .A1(n118), .A2(n74), .ZN(ab_19__2_) );
  NOR2V0P5_8TH40 U873 ( .A1(n117), .A2(n74), .ZN(ab_19__29_) );
  NOR2V0P5_8TH40 U874 ( .A1(n116), .A2(n74), .ZN(ab_19__28_) );
  NOR2V0P5_8TH40 U875 ( .A1(n115), .A2(n74), .ZN(ab_19__27_) );
  NOR2V0P5_8TH40 U876 ( .A1(n114), .A2(n74), .ZN(ab_19__26_) );
  NOR2V0P5_8TH40 U877 ( .A1(n113), .A2(n74), .ZN(ab_19__25_) );
  NOR2V0P5_8TH40 U878 ( .A1(n112), .A2(n74), .ZN(ab_19__24_) );
  NOR2V0P5_8TH40 U879 ( .A1(n111), .A2(n74), .ZN(ab_19__23_) );
  NOR2V0P5_8TH40 U880 ( .A1(n110), .A2(n74), .ZN(ab_19__22_) );
  NOR2V0P5_8TH40 U881 ( .A1(n109), .A2(n74), .ZN(ab_19__21_) );
  NOR2V0P5_8TH40 U882 ( .A1(n108), .A2(n74), .ZN(ab_19__20_) );
  NOR2V0P5_8TH40 U883 ( .A1(n107), .A2(n74), .ZN(ab_19__1_) );
  NOR2V0P5_8TH40 U884 ( .A1(n106), .A2(n74), .ZN(ab_19__19_) );
  NOR2V0P5_8TH40 U885 ( .A1(n105), .A2(n74), .ZN(ab_19__18_) );
  NOR2V0P5_8TH40 U886 ( .A1(n104), .A2(n74), .ZN(ab_19__17_) );
  NOR2V0P5_8TH40 U887 ( .A1(n103), .A2(n74), .ZN(ab_19__16_) );
  NOR2V0P5_8TH40 U888 ( .A1(n102), .A2(n74), .ZN(ab_19__15_) );
  NOR2V0P5_8TH40 U889 ( .A1(n101), .A2(n74), .ZN(ab_19__14_) );
  NOR2V0P5_8TH40 U890 ( .A1(n100), .A2(n74), .ZN(ab_19__13_) );
  NOR2V0P5_8TH40 U891 ( .A1(n99), .A2(n74), .ZN(ab_19__12_) );
  NOR2V0P5_8TH40 U892 ( .A1(n98), .A2(n74), .ZN(ab_19__11_) );
  NOR2V0P5_8TH40 U893 ( .A1(n97), .A2(n74), .ZN(ab_19__10_) );
  NOR2V0P5_8TH40 U894 ( .A1(n96), .A2(n74), .ZN(ab_19__0_) );
  NOR2V0P5_8TH40 U895 ( .A1(n127), .A2(n73), .ZN(ab_18__9_) );
  NOR2V0P5_8TH40 U896 ( .A1(n126), .A2(n73), .ZN(ab_18__8_) );
  NOR2V0P5_8TH40 U897 ( .A1(n125), .A2(n73), .ZN(ab_18__7_) );
  NOR2V0P5_8TH40 U898 ( .A1(n124), .A2(n73), .ZN(ab_18__6_) );
  NOR2V0P5_8TH40 U899 ( .A1(n123), .A2(n73), .ZN(ab_18__5_) );
  NOR2V0P5_8TH40 U900 ( .A1(n122), .A2(n73), .ZN(ab_18__4_) );
  NOR2V0P5_8TH40 U901 ( .A1(n121), .A2(n73), .ZN(ab_18__3_) );
  NOR2V0P5_8TH40 U902 ( .A1(n120), .A2(n73), .ZN(ab_18__31_) );
  NOR2V0P5_8TH40 U903 ( .A1(n119), .A2(n73), .ZN(ab_18__30_) );
  NOR2V0P5_8TH40 U904 ( .A1(n118), .A2(n73), .ZN(ab_18__2_) );
  NOR2V0P5_8TH40 U905 ( .A1(n117), .A2(n73), .ZN(ab_18__29_) );
  NOR2V0P5_8TH40 U906 ( .A1(n116), .A2(n73), .ZN(ab_18__28_) );
  NOR2V0P5_8TH40 U907 ( .A1(n115), .A2(n73), .ZN(ab_18__27_) );
  NOR2V0P5_8TH40 U908 ( .A1(n114), .A2(n73), .ZN(ab_18__26_) );
  NOR2V0P5_8TH40 U909 ( .A1(n113), .A2(n73), .ZN(ab_18__25_) );
  NOR2V0P5_8TH40 U910 ( .A1(n112), .A2(n73), .ZN(ab_18__24_) );
  NOR2V0P5_8TH40 U911 ( .A1(n111), .A2(n73), .ZN(ab_18__23_) );
  NOR2V0P5_8TH40 U912 ( .A1(n110), .A2(n73), .ZN(ab_18__22_) );
  NOR2V0P5_8TH40 U913 ( .A1(n109), .A2(n73), .ZN(ab_18__21_) );
  NOR2V0P5_8TH40 U914 ( .A1(n108), .A2(n73), .ZN(ab_18__20_) );
  NOR2V0P5_8TH40 U915 ( .A1(n107), .A2(n73), .ZN(ab_18__1_) );
  NOR2V0P5_8TH40 U916 ( .A1(n106), .A2(n73), .ZN(ab_18__19_) );
  NOR2V0P5_8TH40 U917 ( .A1(n105), .A2(n73), .ZN(ab_18__18_) );
  NOR2V0P5_8TH40 U918 ( .A1(n104), .A2(n73), .ZN(ab_18__17_) );
  NOR2V0P5_8TH40 U919 ( .A1(n103), .A2(n73), .ZN(ab_18__16_) );
  NOR2V0P5_8TH40 U920 ( .A1(n102), .A2(n73), .ZN(ab_18__15_) );
  NOR2V0P5_8TH40 U921 ( .A1(n101), .A2(n73), .ZN(ab_18__14_) );
  NOR2V0P5_8TH40 U922 ( .A1(n100), .A2(n73), .ZN(ab_18__13_) );
  NOR2V0P5_8TH40 U923 ( .A1(n99), .A2(n73), .ZN(ab_18__12_) );
  NOR2V0P5_8TH40 U924 ( .A1(n98), .A2(n73), .ZN(ab_18__11_) );
  NOR2V0P5_8TH40 U925 ( .A1(n97), .A2(n73), .ZN(ab_18__10_) );
  NOR2V0P5_8TH40 U926 ( .A1(n96), .A2(n73), .ZN(ab_18__0_) );
  NOR2V0P5_8TH40 U927 ( .A1(n127), .A2(n72), .ZN(ab_17__9_) );
  NOR2V0P5_8TH40 U928 ( .A1(n126), .A2(n72), .ZN(ab_17__8_) );
  NOR2V0P5_8TH40 U929 ( .A1(n125), .A2(n72), .ZN(ab_17__7_) );
  NOR2V0P5_8TH40 U930 ( .A1(n124), .A2(n72), .ZN(ab_17__6_) );
  NOR2V0P5_8TH40 U931 ( .A1(n123), .A2(n72), .ZN(ab_17__5_) );
  NOR2V0P5_8TH40 U932 ( .A1(n122), .A2(n72), .ZN(ab_17__4_) );
  NOR2V0P5_8TH40 U933 ( .A1(n121), .A2(n72), .ZN(ab_17__3_) );
  NOR2V0P5_8TH40 U934 ( .A1(n120), .A2(n72), .ZN(ab_17__31_) );
  NOR2V0P5_8TH40 U935 ( .A1(n119), .A2(n72), .ZN(ab_17__30_) );
  NOR2V0P5_8TH40 U936 ( .A1(n118), .A2(n72), .ZN(ab_17__2_) );
  NOR2V0P5_8TH40 U937 ( .A1(n117), .A2(n72), .ZN(ab_17__29_) );
  NOR2V0P5_8TH40 U938 ( .A1(n116), .A2(n72), .ZN(ab_17__28_) );
  NOR2V0P5_8TH40 U939 ( .A1(n115), .A2(n72), .ZN(ab_17__27_) );
  NOR2V0P5_8TH40 U940 ( .A1(n114), .A2(n72), .ZN(ab_17__26_) );
  NOR2V0P5_8TH40 U941 ( .A1(n113), .A2(n72), .ZN(ab_17__25_) );
  NOR2V0P5_8TH40 U942 ( .A1(n112), .A2(n72), .ZN(ab_17__24_) );
  NOR2V0P5_8TH40 U943 ( .A1(n111), .A2(n72), .ZN(ab_17__23_) );
  NOR2V0P5_8TH40 U944 ( .A1(n110), .A2(n72), .ZN(ab_17__22_) );
  NOR2V0P5_8TH40 U945 ( .A1(n109), .A2(n72), .ZN(ab_17__21_) );
  NOR2V0P5_8TH40 U946 ( .A1(n108), .A2(n72), .ZN(ab_17__20_) );
  NOR2V0P5_8TH40 U947 ( .A1(n107), .A2(n72), .ZN(ab_17__1_) );
  NOR2V0P5_8TH40 U948 ( .A1(n106), .A2(n72), .ZN(ab_17__19_) );
  NOR2V0P5_8TH40 U949 ( .A1(n105), .A2(n72), .ZN(ab_17__18_) );
  NOR2V0P5_8TH40 U950 ( .A1(n104), .A2(n72), .ZN(ab_17__17_) );
  NOR2V0P5_8TH40 U951 ( .A1(n103), .A2(n72), .ZN(ab_17__16_) );
  NOR2V0P5_8TH40 U952 ( .A1(n102), .A2(n72), .ZN(ab_17__15_) );
  NOR2V0P5_8TH40 U953 ( .A1(n101), .A2(n72), .ZN(ab_17__14_) );
  NOR2V0P5_8TH40 U954 ( .A1(n100), .A2(n72), .ZN(ab_17__13_) );
  NOR2V0P5_8TH40 U955 ( .A1(n99), .A2(n72), .ZN(ab_17__12_) );
  NOR2V0P5_8TH40 U956 ( .A1(n98), .A2(n72), .ZN(ab_17__11_) );
  NOR2V0P5_8TH40 U957 ( .A1(n97), .A2(n72), .ZN(ab_17__10_) );
  NOR2V0P5_8TH40 U958 ( .A1(n96), .A2(n72), .ZN(ab_17__0_) );
  NOR2V0P5_8TH40 U959 ( .A1(n127), .A2(n71), .ZN(ab_16__9_) );
  NOR2V0P5_8TH40 U960 ( .A1(n126), .A2(n71), .ZN(ab_16__8_) );
  NOR2V0P5_8TH40 U961 ( .A1(n125), .A2(n71), .ZN(ab_16__7_) );
  NOR2V0P5_8TH40 U962 ( .A1(n124), .A2(n71), .ZN(ab_16__6_) );
  NOR2V0P5_8TH40 U963 ( .A1(n123), .A2(n71), .ZN(ab_16__5_) );
  NOR2V0P5_8TH40 U964 ( .A1(n122), .A2(n71), .ZN(ab_16__4_) );
  NOR2V0P5_8TH40 U965 ( .A1(n121), .A2(n71), .ZN(ab_16__3_) );
  NOR2V0P5_8TH40 U966 ( .A1(n120), .A2(n71), .ZN(ab_16__31_) );
  NOR2V0P5_8TH40 U967 ( .A1(n119), .A2(n71), .ZN(ab_16__30_) );
  NOR2V0P5_8TH40 U968 ( .A1(n118), .A2(n71), .ZN(ab_16__2_) );
  NOR2V0P5_8TH40 U969 ( .A1(n117), .A2(n71), .ZN(ab_16__29_) );
  NOR2V0P5_8TH40 U970 ( .A1(n116), .A2(n71), .ZN(ab_16__28_) );
  NOR2V0P5_8TH40 U971 ( .A1(n115), .A2(n71), .ZN(ab_16__27_) );
  NOR2V0P5_8TH40 U972 ( .A1(n114), .A2(n71), .ZN(ab_16__26_) );
  NOR2V0P5_8TH40 U973 ( .A1(n113), .A2(n71), .ZN(ab_16__25_) );
  NOR2V0P5_8TH40 U974 ( .A1(n112), .A2(n71), .ZN(ab_16__24_) );
  NOR2V0P5_8TH40 U975 ( .A1(n111), .A2(n71), .ZN(ab_16__23_) );
  NOR2V0P5_8TH40 U976 ( .A1(n110), .A2(n71), .ZN(ab_16__22_) );
  NOR2V0P5_8TH40 U977 ( .A1(n109), .A2(n71), .ZN(ab_16__21_) );
  NOR2V0P5_8TH40 U978 ( .A1(n108), .A2(n71), .ZN(ab_16__20_) );
  NOR2V0P5_8TH40 U979 ( .A1(n107), .A2(n71), .ZN(ab_16__1_) );
  NOR2V0P5_8TH40 U980 ( .A1(n106), .A2(n71), .ZN(ab_16__19_) );
  NOR2V0P5_8TH40 U981 ( .A1(n105), .A2(n71), .ZN(ab_16__18_) );
  NOR2V0P5_8TH40 U982 ( .A1(n104), .A2(n71), .ZN(ab_16__17_) );
  NOR2V0P5_8TH40 U983 ( .A1(n103), .A2(n71), .ZN(ab_16__16_) );
  NOR2V0P5_8TH40 U984 ( .A1(n102), .A2(n71), .ZN(ab_16__15_) );
  NOR2V0P5_8TH40 U985 ( .A1(n101), .A2(n71), .ZN(ab_16__14_) );
  NOR2V0P5_8TH40 U986 ( .A1(n100), .A2(n71), .ZN(ab_16__13_) );
  NOR2V0P5_8TH40 U987 ( .A1(n99), .A2(n71), .ZN(ab_16__12_) );
  NOR2V0P5_8TH40 U988 ( .A1(n98), .A2(n71), .ZN(ab_16__11_) );
  NOR2V0P5_8TH40 U989 ( .A1(n97), .A2(n71), .ZN(ab_16__10_) );
  NOR2V0P5_8TH40 U990 ( .A1(n96), .A2(n71), .ZN(ab_16__0_) );
  NOR2V0P5_8TH40 U991 ( .A1(n127), .A2(n70), .ZN(ab_15__9_) );
  NOR2V0P5_8TH40 U992 ( .A1(n126), .A2(n70), .ZN(ab_15__8_) );
  NOR2V0P5_8TH40 U993 ( .A1(n125), .A2(n70), .ZN(ab_15__7_) );
  NOR2V0P5_8TH40 U994 ( .A1(n124), .A2(n70), .ZN(ab_15__6_) );
  NOR2V0P5_8TH40 U995 ( .A1(n123), .A2(n70), .ZN(ab_15__5_) );
  NOR2V0P5_8TH40 U996 ( .A1(n122), .A2(n70), .ZN(ab_15__4_) );
  NOR2V0P5_8TH40 U997 ( .A1(n121), .A2(n70), .ZN(ab_15__3_) );
  NOR2V0P5_8TH40 U998 ( .A1(n120), .A2(n70), .ZN(ab_15__31_) );
  NOR2V0P5_8TH40 U999 ( .A1(n119), .A2(n70), .ZN(ab_15__30_) );
  NOR2V0P5_8TH40 U1000 ( .A1(n118), .A2(n70), .ZN(ab_15__2_) );
  NOR2V0P5_8TH40 U1001 ( .A1(n117), .A2(n70), .ZN(ab_15__29_) );
  NOR2V0P5_8TH40 U1002 ( .A1(n116), .A2(n70), .ZN(ab_15__28_) );
  NOR2V0P5_8TH40 U1003 ( .A1(n115), .A2(n70), .ZN(ab_15__27_) );
  NOR2V0P5_8TH40 U1004 ( .A1(n114), .A2(n70), .ZN(ab_15__26_) );
  NOR2V0P5_8TH40 U1005 ( .A1(n113), .A2(n70), .ZN(ab_15__25_) );
  NOR2V0P5_8TH40 U1006 ( .A1(n112), .A2(n70), .ZN(ab_15__24_) );
  NOR2V0P5_8TH40 U1007 ( .A1(n111), .A2(n70), .ZN(ab_15__23_) );
  NOR2V0P5_8TH40 U1008 ( .A1(n110), .A2(n70), .ZN(ab_15__22_) );
  NOR2V0P5_8TH40 U1009 ( .A1(n109), .A2(n70), .ZN(ab_15__21_) );
  NOR2V0P5_8TH40 U1010 ( .A1(n108), .A2(n70), .ZN(ab_15__20_) );
  NOR2V0P5_8TH40 U1011 ( .A1(n107), .A2(n70), .ZN(ab_15__1_) );
  NOR2V0P5_8TH40 U1012 ( .A1(n106), .A2(n70), .ZN(ab_15__19_) );
  NOR2V0P5_8TH40 U1013 ( .A1(n105), .A2(n70), .ZN(ab_15__18_) );
  NOR2V0P5_8TH40 U1014 ( .A1(n104), .A2(n70), .ZN(ab_15__17_) );
  NOR2V0P5_8TH40 U1015 ( .A1(n103), .A2(n70), .ZN(ab_15__16_) );
  NOR2V0P5_8TH40 U1016 ( .A1(n102), .A2(n70), .ZN(ab_15__15_) );
  NOR2V0P5_8TH40 U1017 ( .A1(n101), .A2(n70), .ZN(ab_15__14_) );
  NOR2V0P5_8TH40 U1018 ( .A1(n100), .A2(n70), .ZN(ab_15__13_) );
  NOR2V0P5_8TH40 U1019 ( .A1(n99), .A2(n70), .ZN(ab_15__12_) );
  NOR2V0P5_8TH40 U1020 ( .A1(n98), .A2(n70), .ZN(ab_15__11_) );
  NOR2V0P5_8TH40 U1021 ( .A1(n97), .A2(n70), .ZN(ab_15__10_) );
  NOR2V0P5_8TH40 U1022 ( .A1(n96), .A2(n70), .ZN(ab_15__0_) );
  NOR2V0P5_8TH40 U1023 ( .A1(n127), .A2(n69), .ZN(ab_14__9_) );
  NOR2V0P5_8TH40 U1024 ( .A1(n126), .A2(n69), .ZN(ab_14__8_) );
  NOR2V0P5_8TH40 U1025 ( .A1(n125), .A2(n69), .ZN(ab_14__7_) );
  NOR2V0P5_8TH40 U1026 ( .A1(n124), .A2(n69), .ZN(ab_14__6_) );
  NOR2V0P5_8TH40 U1027 ( .A1(n123), .A2(n69), .ZN(ab_14__5_) );
  NOR2V0P5_8TH40 U1028 ( .A1(n122), .A2(n69), .ZN(ab_14__4_) );
  NOR2V0P5_8TH40 U1029 ( .A1(n121), .A2(n69), .ZN(ab_14__3_) );
  NOR2V0P5_8TH40 U1030 ( .A1(n120), .A2(n69), .ZN(ab_14__31_) );
  NOR2V0P5_8TH40 U1031 ( .A1(n119), .A2(n69), .ZN(ab_14__30_) );
  NOR2V0P5_8TH40 U1032 ( .A1(n118), .A2(n69), .ZN(ab_14__2_) );
  NOR2V0P5_8TH40 U1033 ( .A1(n117), .A2(n69), .ZN(ab_14__29_) );
  NOR2V0P5_8TH40 U1034 ( .A1(n116), .A2(n69), .ZN(ab_14__28_) );
  NOR2V0P5_8TH40 U1035 ( .A1(n115), .A2(n69), .ZN(ab_14__27_) );
  NOR2V0P5_8TH40 U1036 ( .A1(n114), .A2(n69), .ZN(ab_14__26_) );
  NOR2V0P5_8TH40 U1037 ( .A1(n113), .A2(n69), .ZN(ab_14__25_) );
  NOR2V0P5_8TH40 U1038 ( .A1(n112), .A2(n69), .ZN(ab_14__24_) );
  NOR2V0P5_8TH40 U1039 ( .A1(n111), .A2(n69), .ZN(ab_14__23_) );
  NOR2V0P5_8TH40 U1040 ( .A1(n110), .A2(n69), .ZN(ab_14__22_) );
  NOR2V0P5_8TH40 U1041 ( .A1(n109), .A2(n69), .ZN(ab_14__21_) );
  NOR2V0P5_8TH40 U1042 ( .A1(n108), .A2(n69), .ZN(ab_14__20_) );
  NOR2V0P5_8TH40 U1043 ( .A1(n107), .A2(n69), .ZN(ab_14__1_) );
  NOR2V0P5_8TH40 U1044 ( .A1(n106), .A2(n69), .ZN(ab_14__19_) );
  NOR2V0P5_8TH40 U1045 ( .A1(n105), .A2(n69), .ZN(ab_14__18_) );
  NOR2V0P5_8TH40 U1046 ( .A1(n104), .A2(n69), .ZN(ab_14__17_) );
  NOR2V0P5_8TH40 U1047 ( .A1(n103), .A2(n69), .ZN(ab_14__16_) );
  NOR2V0P5_8TH40 U1048 ( .A1(n102), .A2(n69), .ZN(ab_14__15_) );
  NOR2V0P5_8TH40 U1049 ( .A1(n101), .A2(n69), .ZN(ab_14__14_) );
  NOR2V0P5_8TH40 U1050 ( .A1(n100), .A2(n69), .ZN(ab_14__13_) );
  NOR2V0P5_8TH40 U1051 ( .A1(n99), .A2(n69), .ZN(ab_14__12_) );
  NOR2V0P5_8TH40 U1052 ( .A1(n98), .A2(n69), .ZN(ab_14__11_) );
  NOR2V0P5_8TH40 U1053 ( .A1(n97), .A2(n69), .ZN(ab_14__10_) );
  NOR2V0P5_8TH40 U1054 ( .A1(n96), .A2(n69), .ZN(ab_14__0_) );
  NOR2V0P5_8TH40 U1055 ( .A1(n127), .A2(n68), .ZN(ab_13__9_) );
  NOR2V0P5_8TH40 U1056 ( .A1(n126), .A2(n68), .ZN(ab_13__8_) );
  NOR2V0P5_8TH40 U1057 ( .A1(n125), .A2(n68), .ZN(ab_13__7_) );
  NOR2V0P5_8TH40 U1058 ( .A1(n124), .A2(n68), .ZN(ab_13__6_) );
  NOR2V0P5_8TH40 U1059 ( .A1(n123), .A2(n68), .ZN(ab_13__5_) );
  NOR2V0P5_8TH40 U1060 ( .A1(n122), .A2(n68), .ZN(ab_13__4_) );
  NOR2V0P5_8TH40 U1061 ( .A1(n121), .A2(n68), .ZN(ab_13__3_) );
  NOR2V0P5_8TH40 U1062 ( .A1(n120), .A2(n68), .ZN(ab_13__31_) );
  NOR2V0P5_8TH40 U1063 ( .A1(n119), .A2(n68), .ZN(ab_13__30_) );
  NOR2V0P5_8TH40 U1064 ( .A1(n118), .A2(n68), .ZN(ab_13__2_) );
  NOR2V0P5_8TH40 U1065 ( .A1(n117), .A2(n68), .ZN(ab_13__29_) );
  NOR2V0P5_8TH40 U1066 ( .A1(n116), .A2(n68), .ZN(ab_13__28_) );
  NOR2V0P5_8TH40 U1067 ( .A1(n115), .A2(n68), .ZN(ab_13__27_) );
  NOR2V0P5_8TH40 U1068 ( .A1(n114), .A2(n68), .ZN(ab_13__26_) );
  NOR2V0P5_8TH40 U1069 ( .A1(n113), .A2(n68), .ZN(ab_13__25_) );
  NOR2V0P5_8TH40 U1070 ( .A1(n112), .A2(n68), .ZN(ab_13__24_) );
  NOR2V0P5_8TH40 U1071 ( .A1(n111), .A2(n68), .ZN(ab_13__23_) );
  NOR2V0P5_8TH40 U1072 ( .A1(n110), .A2(n68), .ZN(ab_13__22_) );
  NOR2V0P5_8TH40 U1073 ( .A1(n109), .A2(n68), .ZN(ab_13__21_) );
  NOR2V0P5_8TH40 U1074 ( .A1(n108), .A2(n68), .ZN(ab_13__20_) );
  NOR2V0P5_8TH40 U1075 ( .A1(n107), .A2(n68), .ZN(ab_13__1_) );
  NOR2V0P5_8TH40 U1076 ( .A1(n106), .A2(n68), .ZN(ab_13__19_) );
  NOR2V0P5_8TH40 U1077 ( .A1(n105), .A2(n68), .ZN(ab_13__18_) );
  NOR2V0P5_8TH40 U1078 ( .A1(n104), .A2(n68), .ZN(ab_13__17_) );
  NOR2V0P5_8TH40 U1079 ( .A1(n103), .A2(n68), .ZN(ab_13__16_) );
  NOR2V0P5_8TH40 U1080 ( .A1(n102), .A2(n68), .ZN(ab_13__15_) );
  NOR2V0P5_8TH40 U1081 ( .A1(n101), .A2(n68), .ZN(ab_13__14_) );
  NOR2V0P5_8TH40 U1082 ( .A1(n100), .A2(n68), .ZN(ab_13__13_) );
  NOR2V0P5_8TH40 U1083 ( .A1(n99), .A2(n68), .ZN(ab_13__12_) );
  NOR2V0P5_8TH40 U1084 ( .A1(n98), .A2(n68), .ZN(ab_13__11_) );
  NOR2V0P5_8TH40 U1085 ( .A1(n97), .A2(n68), .ZN(ab_13__10_) );
  NOR2V0P5_8TH40 U1086 ( .A1(n96), .A2(n68), .ZN(ab_13__0_) );
  NOR2V0P5_8TH40 U1087 ( .A1(n127), .A2(n67), .ZN(ab_12__9_) );
  NOR2V0P5_8TH40 U1088 ( .A1(n126), .A2(n67), .ZN(ab_12__8_) );
  NOR2V0P5_8TH40 U1089 ( .A1(n125), .A2(n67), .ZN(ab_12__7_) );
  NOR2V0P5_8TH40 U1090 ( .A1(n124), .A2(n67), .ZN(ab_12__6_) );
  NOR2V0P5_8TH40 U1091 ( .A1(n123), .A2(n67), .ZN(ab_12__5_) );
  NOR2V0P5_8TH40 U1092 ( .A1(n122), .A2(n67), .ZN(ab_12__4_) );
  NOR2V0P5_8TH40 U1093 ( .A1(n121), .A2(n67), .ZN(ab_12__3_) );
  NOR2V0P5_8TH40 U1094 ( .A1(n120), .A2(n67), .ZN(ab_12__31_) );
  NOR2V0P5_8TH40 U1095 ( .A1(n119), .A2(n67), .ZN(ab_12__30_) );
  NOR2V0P5_8TH40 U1096 ( .A1(n118), .A2(n67), .ZN(ab_12__2_) );
  NOR2V0P5_8TH40 U1097 ( .A1(n117), .A2(n67), .ZN(ab_12__29_) );
  NOR2V0P5_8TH40 U1098 ( .A1(n116), .A2(n67), .ZN(ab_12__28_) );
  NOR2V0P5_8TH40 U1099 ( .A1(n115), .A2(n67), .ZN(ab_12__27_) );
  NOR2V0P5_8TH40 U1100 ( .A1(n114), .A2(n67), .ZN(ab_12__26_) );
  NOR2V0P5_8TH40 U1101 ( .A1(n113), .A2(n67), .ZN(ab_12__25_) );
  NOR2V0P5_8TH40 U1102 ( .A1(n112), .A2(n67), .ZN(ab_12__24_) );
  NOR2V0P5_8TH40 U1103 ( .A1(n111), .A2(n67), .ZN(ab_12__23_) );
  NOR2V0P5_8TH40 U1104 ( .A1(n110), .A2(n67), .ZN(ab_12__22_) );
  NOR2V0P5_8TH40 U1105 ( .A1(n109), .A2(n67), .ZN(ab_12__21_) );
  NOR2V0P5_8TH40 U1106 ( .A1(n108), .A2(n67), .ZN(ab_12__20_) );
  NOR2V0P5_8TH40 U1107 ( .A1(n107), .A2(n67), .ZN(ab_12__1_) );
  NOR2V0P5_8TH40 U1108 ( .A1(n106), .A2(n67), .ZN(ab_12__19_) );
  NOR2V0P5_8TH40 U1109 ( .A1(n105), .A2(n67), .ZN(ab_12__18_) );
  NOR2V0P5_8TH40 U1110 ( .A1(n104), .A2(n67), .ZN(ab_12__17_) );
  NOR2V0P5_8TH40 U1111 ( .A1(n103), .A2(n67), .ZN(ab_12__16_) );
  NOR2V0P5_8TH40 U1112 ( .A1(n102), .A2(n67), .ZN(ab_12__15_) );
  NOR2V0P5_8TH40 U1113 ( .A1(n101), .A2(n67), .ZN(ab_12__14_) );
  NOR2V0P5_8TH40 U1114 ( .A1(n100), .A2(n67), .ZN(ab_12__13_) );
  NOR2V0P5_8TH40 U1115 ( .A1(n99), .A2(n67), .ZN(ab_12__12_) );
  NOR2V0P5_8TH40 U1116 ( .A1(n98), .A2(n67), .ZN(ab_12__11_) );
  NOR2V0P5_8TH40 U1117 ( .A1(n97), .A2(n67), .ZN(ab_12__10_) );
  NOR2V0P5_8TH40 U1118 ( .A1(n96), .A2(n67), .ZN(ab_12__0_) );
  NOR2V0P5_8TH40 U1119 ( .A1(n127), .A2(n66), .ZN(ab_11__9_) );
  NOR2V0P5_8TH40 U1120 ( .A1(n126), .A2(n66), .ZN(ab_11__8_) );
  NOR2V0P5_8TH40 U1121 ( .A1(n125), .A2(n66), .ZN(ab_11__7_) );
  NOR2V0P5_8TH40 U1122 ( .A1(n124), .A2(n66), .ZN(ab_11__6_) );
  NOR2V0P5_8TH40 U1123 ( .A1(n123), .A2(n66), .ZN(ab_11__5_) );
  NOR2V0P5_8TH40 U1124 ( .A1(n122), .A2(n66), .ZN(ab_11__4_) );
  NOR2V0P5_8TH40 U1125 ( .A1(n121), .A2(n66), .ZN(ab_11__3_) );
  NOR2V0P5_8TH40 U1126 ( .A1(n120), .A2(n66), .ZN(ab_11__31_) );
  NOR2V0P5_8TH40 U1127 ( .A1(n119), .A2(n66), .ZN(ab_11__30_) );
  NOR2V0P5_8TH40 U1128 ( .A1(n118), .A2(n66), .ZN(ab_11__2_) );
  NOR2V0P5_8TH40 U1129 ( .A1(n117), .A2(n66), .ZN(ab_11__29_) );
  NOR2V0P5_8TH40 U1130 ( .A1(n116), .A2(n66), .ZN(ab_11__28_) );
  NOR2V0P5_8TH40 U1131 ( .A1(n115), .A2(n66), .ZN(ab_11__27_) );
  NOR2V0P5_8TH40 U1132 ( .A1(n114), .A2(n66), .ZN(ab_11__26_) );
  NOR2V0P5_8TH40 U1133 ( .A1(n113), .A2(n66), .ZN(ab_11__25_) );
  NOR2V0P5_8TH40 U1134 ( .A1(n112), .A2(n66), .ZN(ab_11__24_) );
  NOR2V0P5_8TH40 U1135 ( .A1(n111), .A2(n66), .ZN(ab_11__23_) );
  NOR2V0P5_8TH40 U1136 ( .A1(n110), .A2(n66), .ZN(ab_11__22_) );
  NOR2V0P5_8TH40 U1137 ( .A1(n109), .A2(n66), .ZN(ab_11__21_) );
  NOR2V0P5_8TH40 U1138 ( .A1(n108), .A2(n66), .ZN(ab_11__20_) );
  NOR2V0P5_8TH40 U1139 ( .A1(n107), .A2(n66), .ZN(ab_11__1_) );
  NOR2V0P5_8TH40 U1140 ( .A1(n106), .A2(n66), .ZN(ab_11__19_) );
  NOR2V0P5_8TH40 U1141 ( .A1(n105), .A2(n66), .ZN(ab_11__18_) );
  NOR2V0P5_8TH40 U1142 ( .A1(n104), .A2(n66), .ZN(ab_11__17_) );
  NOR2V0P5_8TH40 U1143 ( .A1(n103), .A2(n66), .ZN(ab_11__16_) );
  NOR2V0P5_8TH40 U1144 ( .A1(n102), .A2(n66), .ZN(ab_11__15_) );
  NOR2V0P5_8TH40 U1145 ( .A1(n101), .A2(n66), .ZN(ab_11__14_) );
  NOR2V0P5_8TH40 U1146 ( .A1(n100), .A2(n66), .ZN(ab_11__13_) );
  NOR2V0P5_8TH40 U1147 ( .A1(n99), .A2(n66), .ZN(ab_11__12_) );
  NOR2V0P5_8TH40 U1148 ( .A1(n98), .A2(n66), .ZN(ab_11__11_) );
  NOR2V0P5_8TH40 U1149 ( .A1(n97), .A2(n66), .ZN(ab_11__10_) );
  NOR2V0P5_8TH40 U1150 ( .A1(n96), .A2(n66), .ZN(ab_11__0_) );
  NOR2V0P5_8TH40 U1151 ( .A1(n127), .A2(n65), .ZN(ab_10__9_) );
  NOR2V0P5_8TH40 U1152 ( .A1(n126), .A2(n65), .ZN(ab_10__8_) );
  NOR2V0P5_8TH40 U1153 ( .A1(n125), .A2(n65), .ZN(ab_10__7_) );
  NOR2V0P5_8TH40 U1154 ( .A1(n124), .A2(n65), .ZN(ab_10__6_) );
  NOR2V0P5_8TH40 U1155 ( .A1(n123), .A2(n65), .ZN(ab_10__5_) );
  NOR2V0P5_8TH40 U1156 ( .A1(n122), .A2(n65), .ZN(ab_10__4_) );
  NOR2V0P5_8TH40 U1157 ( .A1(n121), .A2(n65), .ZN(ab_10__3_) );
  NOR2V0P5_8TH40 U1158 ( .A1(n120), .A2(n65), .ZN(ab_10__31_) );
  NOR2V0P5_8TH40 U1159 ( .A1(n119), .A2(n65), .ZN(ab_10__30_) );
  NOR2V0P5_8TH40 U1160 ( .A1(n118), .A2(n65), .ZN(ab_10__2_) );
  NOR2V0P5_8TH40 U1161 ( .A1(n117), .A2(n65), .ZN(ab_10__29_) );
  NOR2V0P5_8TH40 U1162 ( .A1(n116), .A2(n65), .ZN(ab_10__28_) );
  NOR2V0P5_8TH40 U1163 ( .A1(n115), .A2(n65), .ZN(ab_10__27_) );
  NOR2V0P5_8TH40 U1164 ( .A1(n114), .A2(n65), .ZN(ab_10__26_) );
  NOR2V0P5_8TH40 U1165 ( .A1(n113), .A2(n65), .ZN(ab_10__25_) );
  NOR2V0P5_8TH40 U1166 ( .A1(n112), .A2(n65), .ZN(ab_10__24_) );
  NOR2V0P5_8TH40 U1167 ( .A1(n111), .A2(n65), .ZN(ab_10__23_) );
  NOR2V0P5_8TH40 U1168 ( .A1(n110), .A2(n65), .ZN(ab_10__22_) );
  NOR2V0P5_8TH40 U1169 ( .A1(n109), .A2(n65), .ZN(ab_10__21_) );
  NOR2V0P5_8TH40 U1170 ( .A1(n108), .A2(n65), .ZN(ab_10__20_) );
  NOR2V0P5_8TH40 U1171 ( .A1(n107), .A2(n65), .ZN(ab_10__1_) );
  NOR2V0P5_8TH40 U1172 ( .A1(n106), .A2(n65), .ZN(ab_10__19_) );
  NOR2V0P5_8TH40 U1173 ( .A1(n105), .A2(n65), .ZN(ab_10__18_) );
  NOR2V0P5_8TH40 U1174 ( .A1(n104), .A2(n65), .ZN(ab_10__17_) );
  NOR2V0P5_8TH40 U1175 ( .A1(n103), .A2(n65), .ZN(ab_10__16_) );
  NOR2V0P5_8TH40 U1176 ( .A1(n102), .A2(n65), .ZN(ab_10__15_) );
  NOR2V0P5_8TH40 U1177 ( .A1(n101), .A2(n65), .ZN(ab_10__14_) );
  NOR2V0P5_8TH40 U1178 ( .A1(n100), .A2(n65), .ZN(ab_10__13_) );
  NOR2V0P5_8TH40 U1179 ( .A1(n99), .A2(n65), .ZN(ab_10__12_) );
  NOR2V0P5_8TH40 U1180 ( .A1(n98), .A2(n65), .ZN(ab_10__11_) );
  NOR2V0P5_8TH40 U1181 ( .A1(n97), .A2(n65), .ZN(ab_10__10_) );
  NOR2V0P5_8TH40 U1182 ( .A1(n96), .A2(n65), .ZN(ab_10__0_) );
  NOR2V0P5_8TH40 U1183 ( .A1(n127), .A2(n64), .ZN(ab_0__9_) );
  NOR2V0P5_8TH40 U1184 ( .A1(n126), .A2(n64), .ZN(ab_0__8_) );
  NOR2V0P5_8TH40 U1185 ( .A1(n125), .A2(n64), .ZN(ab_0__7_) );
  NOR2V0P5_8TH40 U1186 ( .A1(n124), .A2(n64), .ZN(ab_0__6_) );
  NOR2V0P5_8TH40 U1187 ( .A1(n123), .A2(n64), .ZN(ab_0__5_) );
  NOR2V0P5_8TH40 U1188 ( .A1(n122), .A2(n64), .ZN(ab_0__4_) );
  NOR2V0P5_8TH40 U1189 ( .A1(n121), .A2(n64), .ZN(ab_0__3_) );
  NOR2V0P5_8TH40 U1190 ( .A1(n120), .A2(n64), .ZN(ab_0__31_) );
  NOR2V0P5_8TH40 U1191 ( .A1(n119), .A2(n64), .ZN(ab_0__30_) );
  NOR2V0P5_8TH40 U1192 ( .A1(n118), .A2(n64), .ZN(ab_0__2_) );
  NOR2V0P5_8TH40 U1193 ( .A1(n117), .A2(n64), .ZN(ab_0__29_) );
  NOR2V0P5_8TH40 U1194 ( .A1(n116), .A2(n64), .ZN(ab_0__28_) );
  NOR2V0P5_8TH40 U1195 ( .A1(n115), .A2(n64), .ZN(ab_0__27_) );
  NOR2V0P5_8TH40 U1196 ( .A1(n114), .A2(n64), .ZN(ab_0__26_) );
  NOR2V0P5_8TH40 U1197 ( .A1(n113), .A2(n64), .ZN(ab_0__25_) );
  NOR2V0P5_8TH40 U1198 ( .A1(n112), .A2(n64), .ZN(ab_0__24_) );
  NOR2V0P5_8TH40 U1199 ( .A1(n111), .A2(n64), .ZN(ab_0__23_) );
  NOR2V0P5_8TH40 U1200 ( .A1(n110), .A2(n64), .ZN(ab_0__22_) );
  NOR2V0P5_8TH40 U1201 ( .A1(n109), .A2(n64), .ZN(ab_0__21_) );
  NOR2V0P5_8TH40 U1202 ( .A1(n108), .A2(n64), .ZN(ab_0__20_) );
  NOR2V0P5_8TH40 U1203 ( .A1(n107), .A2(n64), .ZN(ab_0__1_) );
  NOR2V0P5_8TH40 U1204 ( .A1(n106), .A2(n64), .ZN(ab_0__19_) );
  NOR2V0P5_8TH40 U1205 ( .A1(n105), .A2(n64), .ZN(ab_0__18_) );
  NOR2V0P5_8TH40 U1206 ( .A1(n104), .A2(n64), .ZN(ab_0__17_) );
  NOR2V0P5_8TH40 U1207 ( .A1(n103), .A2(n64), .ZN(ab_0__16_) );
  NOR2V0P5_8TH40 U1208 ( .A1(n102), .A2(n64), .ZN(ab_0__15_) );
  NOR2V0P5_8TH40 U1209 ( .A1(n101), .A2(n64), .ZN(ab_0__14_) );
  NOR2V0P5_8TH40 U1210 ( .A1(n100), .A2(n64), .ZN(ab_0__13_) );
  NOR2V0P5_8TH40 U1211 ( .A1(n99), .A2(n64), .ZN(ab_0__12_) );
  NOR2V0P5_8TH40 U1212 ( .A1(n98), .A2(n64), .ZN(ab_0__11_) );
  NOR2V0P5_8TH40 U1213 ( .A1(n97), .A2(n64), .ZN(ab_0__10_) );
  NOR2V0P5_8TH40 U1214 ( .A1(n96), .A2(n64), .ZN(PRODUCT[0]) );
endmodule


module inst_execute_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADH1V2C_8TH40 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADH1V2C_8TH40 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADH1V2C_8TH40 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADH1V2C_8TH40 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADH1V2C_8TH40 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADH1V2C_8TH40 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADH1V2C_8TH40 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADH1V2C_8TH40 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADH1V2C_8TH40 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADH1V2C_8TH40 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADH1V2C_8TH40 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADH1V2C_8TH40 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADH1V2C_8TH40 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADH1V2C_8TH40 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADH1V2C_8TH40 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADH1V2C_8TH40 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADH1V2C_8TH40 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADH1V2C_8TH40 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADH1V2C_8TH40 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADH1V2C_8TH40 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADH1V2C_8TH40 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADH1V2C_8TH40 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADH1V2C_8TH40 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADH1V2C_8TH40 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADH1V2C_8TH40 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADH1V2C_8TH40 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADH1V2C_8TH40 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADH1V2C_8TH40 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADH1V2C_8TH40 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADH1V2C_8TH40 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV2_8TH40 U1 ( .I(A[0]), .ZN(SUM[0]) );
  CLKXOR2V2_8TH40 U2 ( .A1(carry[31]), .A2(A[31]), .Z(SUM[31]) );
endmodule


module inst_execute_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADH1V2C_8TH40 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADH1V2C_8TH40 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADH1V2C_8TH40 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADH1V2C_8TH40 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADH1V2C_8TH40 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADH1V2C_8TH40 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADH1V2C_8TH40 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADH1V2C_8TH40 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADH1V2C_8TH40 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADH1V2C_8TH40 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADH1V2C_8TH40 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADH1V2C_8TH40 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADH1V2C_8TH40 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADH1V2C_8TH40 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADH1V2C_8TH40 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADH1V2C_8TH40 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADH1V2C_8TH40 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADH1V2C_8TH40 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADH1V2C_8TH40 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADH1V2C_8TH40 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADH1V2C_8TH40 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADH1V2C_8TH40 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADH1V2C_8TH40 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADH1V2C_8TH40 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADH1V2C_8TH40 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADH1V2C_8TH40 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADH1V2C_8TH40 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADH1V2C_8TH40 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADH1V2C_8TH40 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADH1V2C_8TH40 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV2_8TH40 U1 ( .I(A[0]), .ZN(SUM[0]) );
  CLKXOR2V2_8TH40 U2 ( .A1(carry[31]), .A2(A[31]), .Z(SUM[31]) );
endmodule


module inst_execute_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:2] carry;

  AD1V2C_8TH40 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  AD1V2C_8TH40 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), 
        .S(SUM[30]) );
  AD1V2C_8TH40 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), 
        .S(SUM[29]) );
  AD1V2C_8TH40 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), 
        .S(SUM[28]) );
  AD1V2C_8TH40 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), 
        .S(SUM[27]) );
  AD1V2C_8TH40 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), 
        .S(SUM[26]) );
  AD1V2C_8TH40 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), 
        .S(SUM[25]) );
  AD1V2C_8TH40 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), 
        .S(SUM[24]) );
  AD1V2C_8TH40 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), 
        .S(SUM[23]) );
  AD1V2C_8TH40 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), 
        .S(SUM[22]) );
  AD1V2C_8TH40 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), 
        .S(SUM[21]) );
  AD1V2C_8TH40 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), 
        .S(SUM[20]) );
  AD1V2C_8TH40 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), 
        .S(SUM[19]) );
  AD1V2C_8TH40 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), 
        .S(SUM[18]) );
  AD1V2C_8TH40 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), 
        .S(SUM[17]) );
  AD1V2C_8TH40 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), 
        .S(SUM[16]) );
  AD1V2C_8TH40 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), 
        .S(SUM[15]) );
  AD1V2C_8TH40 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), 
        .S(SUM[14]) );
  AD1V2C_8TH40 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), 
        .S(SUM[13]) );
  AD1V2C_8TH40 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), 
        .S(SUM[12]) );
  AD1V2C_8TH40 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), 
        .S(SUM[11]) );
  AD1V2C_8TH40 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S(SUM[10]) );
  AD1V2C_8TH40 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  AD1V2C_8TH40 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  AD1V2C_8TH40 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  AD1V2C_8TH40 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  AD1V2C_8TH40 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  AD1V2C_8TH40 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  AD1V2C_8TH40 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  AD1V2C_8TH40 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  AD1V2C_8TH40 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1])
         );
  AND2V2_8TH40 U1 ( .A1(A[0]), .A2(B[0]), .Z(n1) );
  XOR2V2_8TH40 U2 ( .A1(A[0]), .A2(B[0]), .Z(SUM[0]) );
endmodule


module inst_execute_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;
  assign DIFF[0] = B[0];

  XOR2V4_8TH40 U1 ( .A1(B[31]), .A2(n30), .Z(DIFF[31]) );
  NAND2V2_8TH40 U2 ( .A1(n29), .A2(n31), .ZN(n30) );
  AND2V2_8TH40 U3 ( .A1(n61), .A2(n60), .Z(n1) );
  AND2V2_8TH40 U4 ( .A1(n1), .A2(n59), .Z(n2) );
  AND2V2_8TH40 U5 ( .A1(n2), .A2(n58), .Z(n3) );
  AND2V2_8TH40 U6 ( .A1(n3), .A2(n57), .Z(n4) );
  AND2V2_8TH40 U7 ( .A1(n4), .A2(n56), .Z(n5) );
  AND2V2_8TH40 U8 ( .A1(n5), .A2(n55), .Z(n6) );
  AND2V2_8TH40 U9 ( .A1(n6), .A2(n54), .Z(n7) );
  AND2V2_8TH40 U10 ( .A1(n7), .A2(n53), .Z(n8) );
  AND2V2_8TH40 U11 ( .A1(n8), .A2(n52), .Z(n9) );
  AND2V2_8TH40 U12 ( .A1(n9), .A2(n51), .Z(n10) );
  AND2V2_8TH40 U13 ( .A1(n10), .A2(n50), .Z(n11) );
  AND2V2_8TH40 U14 ( .A1(n11), .A2(n49), .Z(n12) );
  AND2V2_8TH40 U15 ( .A1(n12), .A2(n48), .Z(n13) );
  AND2V2_8TH40 U16 ( .A1(n13), .A2(n47), .Z(n14) );
  AND2V2_8TH40 U17 ( .A1(n14), .A2(n46), .Z(n15) );
  AND2V2_8TH40 U18 ( .A1(n15), .A2(n45), .Z(n16) );
  AND2V2_8TH40 U19 ( .A1(n16), .A2(n44), .Z(n17) );
  AND2V2_8TH40 U20 ( .A1(n17), .A2(n43), .Z(n18) );
  AND2V2_8TH40 U21 ( .A1(n18), .A2(n42), .Z(n19) );
  AND2V2_8TH40 U22 ( .A1(n19), .A2(n41), .Z(n20) );
  AND2V2_8TH40 U23 ( .A1(n20), .A2(n40), .Z(n21) );
  AND2V2_8TH40 U24 ( .A1(n21), .A2(n39), .Z(n22) );
  AND2V2_8TH40 U25 ( .A1(n22), .A2(n38), .Z(n23) );
  AND2V2_8TH40 U26 ( .A1(n23), .A2(n37), .Z(n24) );
  AND2V2_8TH40 U27 ( .A1(n24), .A2(n36), .Z(n25) );
  AND2V2_8TH40 U28 ( .A1(n25), .A2(n35), .Z(n26) );
  AND2V2_8TH40 U29 ( .A1(n26), .A2(n34), .Z(n27) );
  AND2V2_8TH40 U30 ( .A1(n27), .A2(n33), .Z(n28) );
  AND2V2_8TH40 U31 ( .A1(n28), .A2(n32), .Z(n29) );
  INV2_8TH40 U32 ( .I(B[17]), .ZN(n44) );
  INV2_8TH40 U33 ( .I(B[27]), .ZN(n34) );
  INV2_8TH40 U34 ( .I(B[12]), .ZN(n49) );
  INV2_8TH40 U35 ( .I(B[29]), .ZN(n32) );
  INV2_8TH40 U36 ( .I(B[19]), .ZN(n42) );
  INV2_8TH40 U37 ( .I(B[5]), .ZN(n56) );
  INV2_8TH40 U38 ( .I(B[7]), .ZN(n54) );
  INV2_8TH40 U39 ( .I(B[9]), .ZN(n52) );
  INV2_8TH40 U40 ( .I(B[11]), .ZN(n50) );
  INV2_8TH40 U41 ( .I(B[23]), .ZN(n38) );
  INV2_8TH40 U42 ( .I(B[25]), .ZN(n36) );
  INV2_8TH40 U43 ( .I(B[15]), .ZN(n46) );
  INV2_8TH40 U44 ( .I(B[13]), .ZN(n48) );
  INV2_8TH40 U45 ( .I(B[18]), .ZN(n43) );
  INV2_8TH40 U46 ( .I(B[8]), .ZN(n53) );
  INV2_8TH40 U47 ( .I(B[10]), .ZN(n51) );
  INV2_8TH40 U48 ( .I(B[24]), .ZN(n37) );
  INV2_8TH40 U49 ( .I(B[26]), .ZN(n35) );
  INV2_8TH40 U50 ( .I(B[4]), .ZN(n57) );
  INV2_8TH40 U51 ( .I(B[6]), .ZN(n55) );
  INV2_8TH40 U52 ( .I(B[0]), .ZN(n61) );
  INV2_8TH40 U53 ( .I(B[1]), .ZN(n60) );
  INV2_8TH40 U54 ( .I(B[3]), .ZN(n58) );
  INV2_8TH40 U55 ( .I(B[16]), .ZN(n45) );
  INV2_8TH40 U56 ( .I(B[28]), .ZN(n33) );
  INV2_8TH40 U57 ( .I(B[14]), .ZN(n47) );
  INV2_8TH40 U58 ( .I(B[20]), .ZN(n41) );
  INV2_8TH40 U59 ( .I(B[22]), .ZN(n39) );
  INV2_8TH40 U60 ( .I(B[2]), .ZN(n59) );
  INV2_8TH40 U61 ( .I(B[21]), .ZN(n40) );
  INV2_8TH40 U62 ( .I(B[30]), .ZN(n31) );
  XOR2V2_8TH40 U63 ( .A1(n29), .A2(n31), .Z(DIFF[30]) );
  XOR2V2_8TH40 U64 ( .A1(n28), .A2(n32), .Z(DIFF[29]) );
  XOR2V2_8TH40 U65 ( .A1(n27), .A2(n33), .Z(DIFF[28]) );
  XOR2V2_8TH40 U66 ( .A1(n26), .A2(n34), .Z(DIFF[27]) );
  XOR2V2_8TH40 U67 ( .A1(n25), .A2(n35), .Z(DIFF[26]) );
  XOR2V2_8TH40 U68 ( .A1(n24), .A2(n36), .Z(DIFF[25]) );
  XOR2V2_8TH40 U69 ( .A1(n23), .A2(n37), .Z(DIFF[24]) );
  XOR2V2_8TH40 U70 ( .A1(n22), .A2(n38), .Z(DIFF[23]) );
  XOR2V2_8TH40 U71 ( .A1(n21), .A2(n39), .Z(DIFF[22]) );
  XOR2V2_8TH40 U72 ( .A1(n20), .A2(n40), .Z(DIFF[21]) );
  XOR2V2_8TH40 U73 ( .A1(n19), .A2(n41), .Z(DIFF[20]) );
  XOR2V2_8TH40 U74 ( .A1(n18), .A2(n42), .Z(DIFF[19]) );
  XOR2V2_8TH40 U75 ( .A1(n17), .A2(n43), .Z(DIFF[18]) );
  XOR2V2_8TH40 U76 ( .A1(n16), .A2(n44), .Z(DIFF[17]) );
  XOR2V2_8TH40 U77 ( .A1(n15), .A2(n45), .Z(DIFF[16]) );
  XOR2V2_8TH40 U78 ( .A1(n14), .A2(n46), .Z(DIFF[15]) );
  XOR2V2_8TH40 U79 ( .A1(n13), .A2(n47), .Z(DIFF[14]) );
  XOR2V2_8TH40 U80 ( .A1(n12), .A2(n48), .Z(DIFF[13]) );
  XOR2V2_8TH40 U81 ( .A1(n11), .A2(n49), .Z(DIFF[12]) );
  XOR2V2_8TH40 U82 ( .A1(n10), .A2(n50), .Z(DIFF[11]) );
  XOR2V2_8TH40 U83 ( .A1(n9), .A2(n51), .Z(DIFF[10]) );
  XOR2V2_8TH40 U84 ( .A1(n8), .A2(n52), .Z(DIFF[9]) );
  XOR2V2_8TH40 U85 ( .A1(n7), .A2(n53), .Z(DIFF[8]) );
  XOR2V2_8TH40 U86 ( .A1(n6), .A2(n54), .Z(DIFF[7]) );
  XOR2V2_8TH40 U87 ( .A1(n5), .A2(n55), .Z(DIFF[6]) );
  XOR2V2_8TH40 U88 ( .A1(n4), .A2(n56), .Z(DIFF[5]) );
  XOR2V2_8TH40 U89 ( .A1(n3), .A2(n57), .Z(DIFF[4]) );
  XOR2V2_8TH40 U90 ( .A1(n2), .A2(n58), .Z(DIFF[3]) );
  XOR2V2_8TH40 U91 ( .A1(n1), .A2(n59), .Z(DIFF[2]) );
  XOR2V2_8TH40 U92 ( .A1(n61), .A2(n60), .Z(DIFF[1]) );
endmodule


module inst_execute_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:2] carry;

  AD1V2C_8TH40 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  AD1V2C_8TH40 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), 
        .S(SUM[30]) );
  AD1V2C_8TH40 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), 
        .S(SUM[29]) );
  AD1V2C_8TH40 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), 
        .S(SUM[28]) );
  AD1V2C_8TH40 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), 
        .S(SUM[27]) );
  AD1V2C_8TH40 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), 
        .S(SUM[26]) );
  AD1V2C_8TH40 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), 
        .S(SUM[25]) );
  AD1V2C_8TH40 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), 
        .S(SUM[24]) );
  AD1V2C_8TH40 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), 
        .S(SUM[23]) );
  AD1V2C_8TH40 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), 
        .S(SUM[22]) );
  AD1V2C_8TH40 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), 
        .S(SUM[21]) );
  AD1V2C_8TH40 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), 
        .S(SUM[20]) );
  AD1V2C_8TH40 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), 
        .S(SUM[19]) );
  AD1V2C_8TH40 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), 
        .S(SUM[18]) );
  AD1V2C_8TH40 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), 
        .S(SUM[17]) );
  AD1V2C_8TH40 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), 
        .S(SUM[16]) );
  AD1V2C_8TH40 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), 
        .S(SUM[15]) );
  AD1V2C_8TH40 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), 
        .S(SUM[14]) );
  AD1V2C_8TH40 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), 
        .S(SUM[13]) );
  AD1V2C_8TH40 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), 
        .S(SUM[12]) );
  AD1V2C_8TH40 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), 
        .S(SUM[11]) );
  AD1V2C_8TH40 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S(SUM[10]) );
  AD1V2C_8TH40 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  AD1V2C_8TH40 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  AD1V2C_8TH40 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  AD1V2C_8TH40 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  AD1V2C_8TH40 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  AD1V2C_8TH40 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  AD1V2C_8TH40 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  AD1V2C_8TH40 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  AD1V2C_8TH40 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1])
         );
  AND2V2_8TH40 U1 ( .A1(A[0]), .A2(B[0]), .Z(n1) );
  XOR2V2_8TH40 U2 ( .A1(A[0]), .A2(B[0]), .Z(SUM[0]) );
endmodule


module inst_execute_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159;

  OAI221V2_8TH40 U3 ( .A1(n15), .A2(n1), .B1(n53), .B2(n4), .C(n54), .ZN(B[9])
         );
  OAI221V2_8TH40 U4 ( .A1(n10), .A2(n1), .B1(n58), .B2(n4), .C(n59), .ZN(B[8])
         );
  OAI221V2_8TH40 U5 ( .A1(n11), .A2(n1), .B1(n94), .B2(n4), .C(n142), .ZN(
        B[10]) );
  OAI211V2_8TH40 U6 ( .A1(n13), .A2(n134), .B(n135), .C(n136), .ZN(B[11]) );
  OAI221V2_8TH40 U7 ( .A1(n66), .A2(n1), .B1(n67), .B2(n4), .C(n68), .ZN(B[6])
         );
  OAI221V2_8TH40 U8 ( .A1(n114), .A2(n77), .B1(n109), .B2(n1), .C(n122), .ZN(
        B[13]) );
  OAI221V2_8TH40 U9 ( .A1(n74), .A2(n77), .B1(n115), .B2(n4), .C(n148), .ZN(
        B[0]) );
  AOI222V2_8TH40 U10 ( .A1(n2), .A2(n9), .B1(n80), .B2(n149), .C1(n55), .C2(
        n61), .ZN(n148) );
  OAI221V2_8TH40 U11 ( .A1(n130), .A2(n50), .B1(n124), .B2(n51), .C(n152), 
        .ZN(n149) );
  OAI221V2_8TH40 U12 ( .A1(n62), .A2(n77), .B1(n78), .B2(n4), .C(n79), .ZN(
        B[3]) );
  AOI222V2_8TH40 U13 ( .A1(n2), .A2(n21), .B1(n80), .B2(n81), .C1(n55), .C2(
        n65), .ZN(n79) );
  OAI221V2_8TH40 U14 ( .A1(n25), .A2(n49), .B1(n24), .B2(n50), .C(n82), .ZN(
        n81) );
  AOI221V2_8TH40 U15 ( .A1(n56), .A2(n97), .B1(n22), .B2(n96), .C(n113), .ZN(
        n104) );
  AOI221V2_8TH40 U16 ( .A1(n103), .A2(n97), .B1(n70), .B2(n96), .C(n111), .ZN(
        n86) );
  AOI221V2_8TH40 U17 ( .A1(n60), .A2(n97), .B1(n17), .B2(n96), .C(n154), .ZN(
        n115) );
  OAI221V2_8TH40 U18 ( .A1(n71), .A2(n77), .B1(n104), .B2(n4), .C(n105), .ZN(
        B[1]) );
  AOI222V2_8TH40 U19 ( .A1(n2), .A2(n14), .B1(n80), .B2(n106), .C1(n55), .C2(
        n57), .ZN(n105) );
  OAI221V2_8TH40 U20 ( .A1(n25), .A2(n51), .B1(n24), .B2(n52), .C(n108), .ZN(
        n106) );
  OAI221V2_8TH40 U21 ( .A1(n66), .A2(n77), .B1(n86), .B2(n4), .C(n87), .ZN(
        B[2]) );
  AOI222V2_8TH40 U22 ( .A1(n2), .A2(n12), .B1(n80), .B2(n88), .C1(n55), .C2(
        n69), .ZN(n87) );
  OAI221V2_8TH40 U23 ( .A1(n25), .A2(n50), .B1(n24), .B2(n51), .C(n89), .ZN(
        n88) );
  OAI221V2_8TH40 U24 ( .A1(n116), .A2(n77), .B1(n117), .B2(n1), .C(n118), .ZN(
        B[15]) );
  OAI221V2_8TH40 U25 ( .A1(n131), .A2(n77), .B1(n132), .B2(n1), .C(n133), .ZN(
        B[12]) );
  OAI221V2_8TH40 U26 ( .A1(n62), .A2(n1), .B1(n63), .B2(n4), .C(n64), .ZN(B[7]) );
  OAI221V2_8TH40 U27 ( .A1(n71), .A2(n1), .B1(n72), .B2(n4), .C(n73), .ZN(B[5]) );
  OAI221V2_8TH40 U28 ( .A1(n74), .A2(n1), .B1(n75), .B2(n4), .C(n76), .ZN(B[4]) );
  OAI221V2_8TH40 U29 ( .A1(n130), .A2(n36), .B1(n37), .B2(n124), .C(n144), 
        .ZN(n70) );
  OAI221V2_8TH40 U30 ( .A1(n25), .A2(n33), .B1(n24), .B2(n34), .C(n141), .ZN(
        n101) );
  AOI221V2_8TH40 U31 ( .A1(n126), .A2(A[29]), .B1(n127), .B2(A[28]), .C(n156), 
        .ZN(n92) );
  AOI221V2_8TH40 U32 ( .A1(n126), .A2(A[14]), .B1(n127), .B2(A[13]), .C(n128), 
        .ZN(n109) );
  AOI221V2_8TH40 U33 ( .A1(n126), .A2(A[15]), .B1(n127), .B2(A[14]), .C(n145), 
        .ZN(n120) );
  AOI221V2_8TH40 U34 ( .A1(n126), .A2(A[13]), .B1(n127), .B2(A[12]), .C(n153), 
        .ZN(n132) );
  OAI22V2_8TH40 U35 ( .A1(n39), .A2(n130), .B1(n40), .B2(n124), .ZN(n138) );
  AOI221V2_8TH40 U36 ( .A1(A[20]), .A2(n126), .B1(A[19]), .B2(n127), .C(n139), 
        .ZN(n116) );
  AOI221V2_8TH40 U37 ( .A1(n126), .A2(A[18]), .B1(n127), .B2(A[17]), .C(n129), 
        .ZN(n114) );
  AOI221V2_8TH40 U38 ( .A1(n126), .A2(A[17]), .B1(n127), .B2(A[16]), .C(n157), 
        .ZN(n131) );
  OAI221V2_8TH40 U39 ( .A1(n25), .A2(n35), .B1(n24), .B2(n36), .C(n123), .ZN(
        n56) );
  OAI221V2_8TH40 U40 ( .A1(n25), .A2(n36), .B1(n37), .B2(n24), .C(n158), .ZN(
        n60) );
  OAI221V2_8TH40 U41 ( .A1(n25), .A2(n34), .B1(n24), .B2(n35), .C(n143), .ZN(
        n103) );
  OAI221V2_8TH40 U42 ( .A1(n25), .A2(n31), .B1(n24), .B2(n32), .C(n125), .ZN(
        n95) );
  OAI221V2_8TH40 U43 ( .A1(n25), .A2(n32), .B1(n24), .B2(n33), .C(n155), .ZN(
        n98) );
  OAI221V2_8TH40 U44 ( .A1(n25), .A2(n42), .B1(n24), .B2(n43), .C(n147), .ZN(
        n69) );
  OAI221V2_8TH40 U45 ( .A1(n25), .A2(n44), .B1(n24), .B2(n45), .C(n150), .ZN(
        n61) );
  OAI221V2_8TH40 U46 ( .A1(n25), .A2(n43), .B1(n24), .B2(n44), .C(n107), .ZN(
        n57) );
  AO221V2_8TH40 U47 ( .A1(n126), .A2(A[28]), .B1(n127), .B2(A[27]), .C(n140), 
        .Z(n99) );
  OA221V2_8TH40 U48 ( .A1(n25), .A2(n46), .B1(n24), .B2(n47), .C(n90), .Z(n66)
         );
  OA221V2_8TH40 U49 ( .A1(n25), .A2(n47), .B1(n24), .B2(n48), .C(n110), .Z(n71) );
  OA221V2_8TH40 U50 ( .A1(n25), .A2(n45), .B1(n24), .B2(n46), .C(n83), .Z(n62)
         );
  OA221V2_8TH40 U51 ( .A1(n25), .A2(n48), .B1(n24), .B2(n49), .C(n159), .Z(n74) );
  INV2_8TH40 U52 ( .I(n77), .ZN(n3) );
  INV2_8TH40 U53 ( .I(n93), .ZN(n7) );
  INV2_8TH40 U54 ( .I(n61), .ZN(n10) );
  INV2_8TH40 U55 ( .I(n57), .ZN(n15) );
  INV2_8TH40 U56 ( .I(n69), .ZN(n11) );
  INV2_8TH40 U57 ( .I(n127), .ZN(n24) );
  INV2_8TH40 U58 ( .I(n126), .ZN(n25) );
  INV2_8TH40 U59 ( .I(n70), .ZN(n19) );
  INV2_8TH40 U60 ( .I(n80), .ZN(n1) );
  INV2_8TH40 U61 ( .I(n124), .ZN(n16) );
  INV2_8TH40 U62 ( .I(n130), .ZN(n23) );
  INV2_8TH40 U63 ( .I(n96), .ZN(n6) );
  INV2_8TH40 U64 ( .I(n92), .ZN(n18) );
  INV2_8TH40 U65 ( .I(n134), .ZN(n2) );
  INV2_8TH40 U66 ( .I(n132), .ZN(n9) );
  INV2_8TH40 U67 ( .I(n109), .ZN(n14) );
  INV2_8TH40 U68 ( .I(n120), .ZN(n12) );
  INV2_8TH40 U69 ( .I(n117), .ZN(n21) );
  INV2_8TH40 U70 ( .I(n114), .ZN(n22) );
  INV2_8TH40 U71 ( .I(n131), .ZN(n17) );
  INV2_8TH40 U72 ( .I(n116), .ZN(n20) );
  INV2_8TH40 U73 ( .I(n101), .ZN(n13) );
  INV2_8TH40 U74 ( .I(A[17]), .ZN(n40) );
  INV2_8TH40 U75 ( .I(A[27]), .ZN(n30) );
  INV2_8TH40 U76 ( .I(A[12]), .ZN(n41) );
  INV2_8TH40 U77 ( .I(SH[4]), .ZN(n4) );
  INV2_8TH40 U78 ( .I(SH[2]), .ZN(n8) );
  INV2_8TH40 U79 ( .I(SH[3]), .ZN(n5) );
  INV2_8TH40 U80 ( .I(SH[0]), .ZN(n26) );
  INV2_8TH40 U81 ( .I(A[31]), .ZN(n27) );
  INV2_8TH40 U82 ( .I(A[21]), .ZN(n36) );
  INV2_8TH40 U83 ( .I(A[30]), .ZN(n28) );
  INV2_8TH40 U84 ( .I(A[3]), .ZN(n50) );
  INV2_8TH40 U85 ( .I(A[22]), .ZN(n35) );
  INV2_8TH40 U86 ( .I(A[20]), .ZN(n37) );
  INV2_8TH40 U87 ( .I(A[2]), .ZN(n51) );
  INV2_8TH40 U88 ( .I(A[5]), .ZN(n48) );
  INV2_8TH40 U89 ( .I(A[7]), .ZN(n46) );
  INV2_8TH40 U90 ( .I(A[9]), .ZN(n44) );
  INV2_8TH40 U91 ( .I(A[11]), .ZN(n42) );
  INV2_8TH40 U92 ( .I(A[23]), .ZN(n34) );
  INV2_8TH40 U93 ( .I(A[25]), .ZN(n32) );
  INV2_8TH40 U94 ( .I(A[29]), .ZN(n29) );
  INV2_8TH40 U95 ( .I(A[19]), .ZN(n38) );
  INV2_8TH40 U96 ( .I(A[8]), .ZN(n45) );
  INV2_8TH40 U97 ( .I(A[10]), .ZN(n43) );
  INV2_8TH40 U98 ( .I(A[24]), .ZN(n33) );
  INV2_8TH40 U99 ( .I(A[26]), .ZN(n31) );
  INV2_8TH40 U100 ( .I(A[6]), .ZN(n47) );
  INV2_8TH40 U101 ( .I(A[4]), .ZN(n49) );
  INV2_8TH40 U102 ( .I(A[18]), .ZN(n39) );
  INV2_8TH40 U103 ( .I(A[1]), .ZN(n52) );
  AOI222V0_8TH40 U104 ( .A1(n3), .A2(n14), .B1(n55), .B2(n22), .C1(n2), .C2(
        n56), .ZN(n54) );
  AOI222V0_8TH40 U105 ( .A1(n3), .A2(n9), .B1(n55), .B2(n17), .C1(n2), .C2(n60), .ZN(n59) );
  AOI222V0_8TH40 U106 ( .A1(n3), .A2(n65), .B1(n55), .B2(n21), .C1(n2), .C2(
        n20), .ZN(n64) );
  AOI222V0_8TH40 U107 ( .A1(n3), .A2(n69), .B1(n55), .B2(n12), .C1(n2), .C2(
        n70), .ZN(n68) );
  AOI222V0_8TH40 U108 ( .A1(n3), .A2(n57), .B1(n55), .B2(n14), .C1(n2), .C2(
        n22), .ZN(n73) );
  AOI222V0_8TH40 U109 ( .A1(n3), .A2(n61), .B1(n55), .B2(n9), .C1(n2), .C2(n17), .ZN(n76) );
  AOI22V0_8TH40 U110 ( .A1(A[6]), .A2(n23), .B1(A[5]), .B2(n16), .ZN(n82) );
  AOI22V0_8TH40 U111 ( .A1(A[10]), .A2(n23), .B1(A[9]), .B2(n16), .ZN(n83) );
  AND2V0_8TH40 U112 ( .A1(n84), .A2(n80), .Z(B[31]) );
  INOR2V0_8TH40 U113 ( .A1(n85), .B1(n1), .ZN(B[30]) );
  AOI22V0_8TH40 U114 ( .A1(A[5]), .A2(n23), .B1(A[4]), .B2(n16), .ZN(n89) );
  AOI22V0_8TH40 U115 ( .A1(A[9]), .A2(n23), .B1(A[8]), .B2(n16), .ZN(n90) );
  AND2V0_8TH40 U116 ( .A1(n91), .A2(n80), .Z(B[29]) );
  NOR2V0P5_8TH40 U117 ( .A1(n92), .A2(n1), .ZN(B[28]) );
  NOR3V0P5_8TH40 U118 ( .A1(n93), .A2(SH[4]), .A3(SH[3]), .ZN(B[27]) );
  NOR2V0P5_8TH40 U119 ( .A1(SH[4]), .A2(n94), .ZN(B[26]) );
  NOR2V0P5_8TH40 U120 ( .A1(SH[4]), .A2(n53), .ZN(B[25]) );
  AOI22V0_8TH40 U121 ( .A1(n95), .A2(n96), .B1(n91), .B2(n97), .ZN(n53) );
  NOR2V0P5_8TH40 U122 ( .A1(SH[4]), .A2(n58), .ZN(B[24]) );
  AOI22V0_8TH40 U123 ( .A1(n98), .A2(n96), .B1(n18), .B2(n97), .ZN(n58) );
  NOR2V0P5_8TH40 U124 ( .A1(SH[4]), .A2(n63), .ZN(B[23]) );
  AOI222V0_8TH40 U125 ( .A1(n99), .A2(n97), .B1(n84), .B2(n100), .C1(n101), 
        .C2(n96), .ZN(n63) );
  NOR2V0P5_8TH40 U126 ( .A1(SH[4]), .A2(n67), .ZN(B[22]) );
  AOI222V0_8TH40 U127 ( .A1(n102), .A2(n97), .B1(n85), .B2(n100), .C1(n103), 
        .C2(n96), .ZN(n67) );
  NOR2V0P5_8TH40 U128 ( .A1(SH[4]), .A2(n72), .ZN(B[21]) );
  AOI222V0_8TH40 U129 ( .A1(n95), .A2(n97), .B1(n91), .B2(n100), .C1(n56), 
        .C2(n96), .ZN(n72) );
  NOR2V0P5_8TH40 U130 ( .A1(SH[4]), .A2(n75), .ZN(B[20]) );
  AOI222V0_8TH40 U131 ( .A1(n98), .A2(n97), .B1(n18), .B2(n100), .C1(n60), 
        .C2(n96), .ZN(n75) );
  AOI22V0_8TH40 U132 ( .A1(A[12]), .A2(n23), .B1(A[11]), .B2(n16), .ZN(n107)
         );
  AOI22V0_8TH40 U133 ( .A1(A[4]), .A2(n23), .B1(A[3]), .B2(n16), .ZN(n108) );
  AOI22V0_8TH40 U134 ( .A1(A[8]), .A2(n23), .B1(A[7]), .B2(n16), .ZN(n110) );
  NOR2V0P5_8TH40 U135 ( .A1(SH[4]), .A2(n78), .ZN(B[19]) );
  AOI222V0_8TH40 U136 ( .A1(n20), .A2(n96), .B1(n101), .B2(n97), .C1(n7), .C2(
        SH[3]), .ZN(n78) );
  NOR2V0P5_8TH40 U137 ( .A1(SH[4]), .A2(n86), .ZN(B[18]) );
  AO22V0_8TH40 U138 ( .A1(n112), .A2(n85), .B1(n100), .B2(n102), .Z(n111) );
  NOR2V0P5_8TH40 U139 ( .A1(SH[4]), .A2(n104), .ZN(B[17]) );
  AO22V0_8TH40 U140 ( .A1(n112), .A2(n91), .B1(n100), .B2(n95), .Z(n113) );
  NOR2V0P5_8TH40 U141 ( .A1(SH[4]), .A2(n115), .ZN(B[16]) );
  AOI222V0_8TH40 U142 ( .A1(n2), .A2(n99), .B1(n119), .B2(n84), .C1(n55), .C2(
        n101), .ZN(n118) );
  OAI221V0_8TH40 U143 ( .A1(n19), .A2(n77), .B1(n120), .B2(n1), .C(n121), .ZN(
        B[14]) );
  AOI222V0_8TH40 U144 ( .A1(n2), .A2(n102), .B1(n119), .B2(n85), .C1(n55), 
        .C2(n103), .ZN(n121) );
  AOI222V0_8TH40 U145 ( .A1(n2), .A2(n95), .B1(n119), .B2(n91), .C1(n55), .C2(
        n56), .ZN(n122) );
  AOI22V0_8TH40 U146 ( .A1(A[24]), .A2(n23), .B1(A[23]), .B2(n16), .ZN(n123)
         );
  OAI222V0_8TH40 U147 ( .A1(n25), .A2(n28), .B1(n124), .B2(n27), .C1(n24), 
        .C2(n29), .ZN(n91) );
  AOI22V0_8TH40 U148 ( .A1(A[28]), .A2(n23), .B1(A[27]), .B2(n16), .ZN(n125)
         );
  AO22V0_8TH40 U149 ( .A1(A[16]), .A2(n23), .B1(A[15]), .B2(n16), .Z(n128) );
  OAI22V0_8TH40 U150 ( .A1(n37), .A2(n130), .B1(n38), .B2(n124), .ZN(n129) );
  AOI222V0_8TH40 U151 ( .A1(n2), .A2(n98), .B1(n119), .B2(n18), .C1(n55), .C2(
        n60), .ZN(n133) );
  NOR2V0P5_8TH40 U152 ( .A1(n4), .A2(n6), .ZN(n119) );
  AOI22V0_8TH40 U153 ( .A1(n3), .A2(n21), .B1(n80), .B2(n65), .ZN(n136) );
  OAI221V0_8TH40 U154 ( .A1(n25), .A2(n41), .B1(n24), .B2(n42), .C(n137), .ZN(
        n65) );
  AOI22V0_8TH40 U155 ( .A1(A[14]), .A2(n23), .B1(A[13]), .B2(n16), .ZN(n137)
         );
  AOI221V0_8TH40 U156 ( .A1(n126), .A2(A[16]), .B1(n127), .B2(A[15]), .C(n138), 
        .ZN(n117) );
  AOI32V0_8TH40 U157 ( .A1(n7), .A2(n5), .A3(SH[4]), .B1(n55), .B2(n20), .ZN(
        n135) );
  OAI22V0_8TH40 U158 ( .A1(n35), .A2(n130), .B1(n36), .B2(n124), .ZN(n139) );
  MUX2NV0_8TH40 U159 ( .I0(n84), .I1(n99), .S(n8), .ZN(n93) );
  OAI22V0_8TH40 U160 ( .A1(n28), .A2(n130), .B1(n29), .B2(n124), .ZN(n140) );
  NOR2V0P5_8TH40 U161 ( .A1(n27), .A2(n24), .ZN(n84) );
  AOI22V0_8TH40 U162 ( .A1(A[26]), .A2(n23), .B1(A[25]), .B2(n16), .ZN(n141)
         );
  AOI222V0_8TH40 U163 ( .A1(n3), .A2(n12), .B1(n55), .B2(n70), .C1(n2), .C2(
        n103), .ZN(n142) );
  AOI22V0_8TH40 U164 ( .A1(A[25]), .A2(n23), .B1(A[24]), .B2(n16), .ZN(n143)
         );
  AOI22V0_8TH40 U165 ( .A1(n126), .A2(A[19]), .B1(n127), .B2(A[18]), .ZN(n144)
         );
  AO22V0_8TH40 U166 ( .A1(A[17]), .A2(n23), .B1(A[16]), .B2(n16), .Z(n145) );
  AOI22V0_8TH40 U167 ( .A1(n102), .A2(n96), .B1(n85), .B2(n97), .ZN(n94) );
  OAI22V0_8TH40 U168 ( .A1(n24), .A2(n28), .B1(n25), .B2(n27), .ZN(n85) );
  OAI221V0_8TH40 U169 ( .A1(n25), .A2(n30), .B1(n24), .B2(n31), .C(n146), .ZN(
        n102) );
  AOI22V0_8TH40 U170 ( .A1(A[29]), .A2(n23), .B1(A[28]), .B2(n16), .ZN(n146)
         );
  AOI22V0_8TH40 U171 ( .A1(A[13]), .A2(n23), .B1(A[12]), .B2(n16), .ZN(n147)
         );
  AOI22V0_8TH40 U172 ( .A1(A[11]), .A2(n23), .B1(A[10]), .B2(n16), .ZN(n150)
         );
  AND2V0_8TH40 U173 ( .A1(n151), .A2(n8), .Z(n55) );
  AOI22V0_8TH40 U174 ( .A1(A[1]), .A2(n126), .B1(A[0]), .B2(n127), .ZN(n152)
         );
  NOR2V0P5_8TH40 U175 ( .A1(n6), .A2(SH[4]), .ZN(n80) );
  AO22V0_8TH40 U176 ( .A1(A[15]), .A2(n23), .B1(A[14]), .B2(n16), .Z(n153) );
  CLKNAND2V1_8TH40 U177 ( .A1(SH[2]), .A2(n151), .ZN(n134) );
  NOR2V0P5_8TH40 U178 ( .A1(n5), .A2(SH[4]), .ZN(n151) );
  AO22V0_8TH40 U179 ( .A1(n112), .A2(n18), .B1(n100), .B2(n98), .Z(n154) );
  AOI22V0_8TH40 U180 ( .A1(A[27]), .A2(n23), .B1(A[26]), .B2(n16), .ZN(n155)
         );
  NOR2V0P5_8TH40 U181 ( .A1(n5), .A2(SH[2]), .ZN(n100) );
  OAI22V0_8TH40 U182 ( .A1(n27), .A2(n130), .B1(n28), .B2(n124), .ZN(n156) );
  NOR2V0P5_8TH40 U183 ( .A1(n8), .A2(n5), .ZN(n112) );
  NOR2V0P5_8TH40 U184 ( .A1(SH[2]), .A2(SH[3]), .ZN(n96) );
  OAI22V0_8TH40 U185 ( .A1(n38), .A2(n130), .B1(n39), .B2(n124), .ZN(n157) );
  AOI22V0_8TH40 U186 ( .A1(A[23]), .A2(n23), .B1(A[22]), .B2(n16), .ZN(n158)
         );
  CLKNAND2V1_8TH40 U187 ( .A1(n97), .A2(n4), .ZN(n77) );
  NOR2V0P5_8TH40 U188 ( .A1(n8), .A2(SH[3]), .ZN(n97) );
  AOI22V0_8TH40 U189 ( .A1(A[7]), .A2(n23), .B1(A[6]), .B2(n16), .ZN(n159) );
  CLKNAND2V1_8TH40 U190 ( .A1(SH[1]), .A2(n26), .ZN(n124) );
  CLKNAND2V1_8TH40 U191 ( .A1(SH[1]), .A2(SH[0]), .ZN(n130) );
  NOR2V0P5_8TH40 U192 ( .A1(SH[0]), .A2(SH[1]), .ZN(n127) );
  NOR2V0P5_8TH40 U193 ( .A1(n26), .A2(SH[1]), .ZN(n126) );
endmodule


module inst_execute_DW01_add_3 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:2] carry;

  AD1V2C_8TH40 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .S(SUM[63]) );
  AD1V2C_8TH40 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), 
        .S(SUM[62]) );
  AD1V2C_8TH40 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), 
        .S(SUM[61]) );
  AD1V2C_8TH40 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), 
        .S(SUM[60]) );
  AD1V2C_8TH40 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), 
        .S(SUM[59]) );
  AD1V2C_8TH40 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), 
        .S(SUM[58]) );
  AD1V2C_8TH40 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), 
        .S(SUM[57]) );
  AD1V2C_8TH40 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), 
        .S(SUM[56]) );
  AD1V2C_8TH40 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), 
        .S(SUM[55]) );
  AD1V2C_8TH40 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), 
        .S(SUM[54]) );
  AD1V2C_8TH40 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), 
        .S(SUM[53]) );
  AD1V2C_8TH40 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), 
        .S(SUM[52]) );
  AD1V2C_8TH40 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), 
        .S(SUM[51]) );
  AD1V2C_8TH40 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), 
        .S(SUM[50]) );
  AD1V2C_8TH40 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), 
        .S(SUM[49]) );
  AD1V2C_8TH40 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), 
        .S(SUM[48]) );
  AD1V2C_8TH40 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), 
        .S(SUM[47]) );
  AD1V2C_8TH40 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), 
        .S(SUM[46]) );
  AD1V2C_8TH40 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), 
        .S(SUM[45]) );
  AD1V2C_8TH40 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), 
        .S(SUM[44]) );
  AD1V2C_8TH40 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), 
        .S(SUM[43]) );
  AD1V2C_8TH40 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), 
        .S(SUM[42]) );
  AD1V2C_8TH40 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), 
        .S(SUM[41]) );
  AD1V2C_8TH40 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), 
        .S(SUM[40]) );
  AD1V2C_8TH40 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), 
        .S(SUM[39]) );
  AD1V2C_8TH40 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), 
        .S(SUM[38]) );
  AD1V2C_8TH40 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), 
        .S(SUM[37]) );
  AD1V2C_8TH40 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), 
        .S(SUM[36]) );
  AD1V2C_8TH40 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), 
        .S(SUM[35]) );
  AD1V2C_8TH40 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), 
        .S(SUM[34]) );
  AD1V2C_8TH40 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), 
        .S(SUM[33]) );
  AD1V2C_8TH40 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), 
        .S(SUM[32]) );
  AD1V2C_8TH40 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), 
        .S(SUM[31]) );
  AD1V2C_8TH40 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), 
        .S(SUM[30]) );
  AD1V2C_8TH40 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), 
        .S(SUM[29]) );
  AD1V2C_8TH40 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), 
        .S(SUM[28]) );
  AD1V2C_8TH40 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), 
        .S(SUM[27]) );
  AD1V2C_8TH40 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), 
        .S(SUM[26]) );
  AD1V2C_8TH40 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), 
        .S(SUM[25]) );
  AD1V2C_8TH40 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), 
        .S(SUM[24]) );
  AD1V2C_8TH40 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), 
        .S(SUM[23]) );
  AD1V2C_8TH40 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), 
        .S(SUM[22]) );
  AD1V2C_8TH40 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), 
        .S(SUM[21]) );
  AD1V2C_8TH40 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), 
        .S(SUM[20]) );
  AD1V2C_8TH40 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), 
        .S(SUM[19]) );
  AD1V2C_8TH40 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), 
        .S(SUM[18]) );
  AD1V2C_8TH40 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), 
        .S(SUM[17]) );
  AD1V2C_8TH40 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), 
        .S(SUM[16]) );
  AD1V2C_8TH40 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), 
        .S(SUM[15]) );
  AD1V2C_8TH40 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), 
        .S(SUM[14]) );
  AD1V2C_8TH40 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), 
        .S(SUM[13]) );
  AD1V2C_8TH40 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), 
        .S(SUM[12]) );
  AD1V2C_8TH40 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), 
        .S(SUM[11]) );
  AD1V2C_8TH40 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S(SUM[10]) );
  AD1V2C_8TH40 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  AD1V2C_8TH40 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  AD1V2C_8TH40 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  AD1V2C_8TH40 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  AD1V2C_8TH40 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  AD1V2C_8TH40 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  AD1V2C_8TH40 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  AD1V2C_8TH40 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  AD1V2C_8TH40 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1])
         );
  AND2V2_8TH40 U1 ( .A1(A[0]), .A2(B[0]), .Z(n1) );
  XOR2V2_8TH40 U2 ( .A1(A[0]), .A2(B[0]), .Z(SUM[0]) );
endmodule


module inst_execute_DW01_cmp6_2 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105;

  AOI32V2_8TH40 U1 ( .A1(n49), .A2(n50), .A3(n78), .B1(B[24]), .B2(n4), .ZN(
        n77) );
  AOI32V2_8TH40 U2 ( .A1(n55), .A2(n56), .A3(n84), .B1(B[18]), .B2(n7), .ZN(
        n83) );
  AOI32V2_8TH40 U3 ( .A1(n63), .A2(n64), .A3(n90), .B1(B[12]), .B2(n10), .ZN(
        n89) );
  OAI211V2_8TH40 U4 ( .A1(n104), .A2(n15), .B(n105), .C(n68), .ZN(n103) );
  OAI21V2_8TH40 U5 ( .A1(A[27]), .A2(n18), .B(n75), .ZN(n74) );
  OAI21V2_8TH40 U6 ( .A1(A[21]), .A2(n21), .B(n81), .ZN(n80) );
  OAI21V2_8TH40 U7 ( .A1(A[15]), .A2(n24), .B(n87), .ZN(n86) );
  OAI21V2_8TH40 U8 ( .A1(A[9]), .A2(n27), .B(n93), .ZN(n92) );
  AOI32V2_8TH40 U9 ( .A1(n42), .A2(n43), .A3(n72), .B1(B[30]), .B2(n1), .ZN(
        n71) );
  NOR4V2_8TH40 U10 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n36) );
  NAND4V2_8TH40 U11 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .ZN(NE) );
  NOR2V2_8TH40 U12 ( .A1(n58), .A2(n59), .ZN(n35) );
  OAI21V2_8TH40 U13 ( .A1(A[29]), .A2(n17), .B(n73), .ZN(n72) );
  AOI32V2_8TH40 U14 ( .A1(n67), .A2(n94), .A3(n95), .B1(B[8]), .B2(n12), .ZN(
        n93) );
  AOI32V2_8TH40 U15 ( .A1(n61), .A2(n62), .A3(n88), .B1(B[14]), .B2(n9), .ZN(
        n87) );
  AOI32V2_8TH40 U16 ( .A1(n53), .A2(n54), .A3(n82), .B1(B[20]), .B2(n6), .ZN(
        n81) );
  AOI32V2_8TH40 U17 ( .A1(n47), .A2(n48), .A3(n76), .B1(B[26]), .B2(n3), .ZN(
        n75) );
  OAI21V2_8TH40 U18 ( .A1(A[7]), .A2(n28), .B(n96), .ZN(n95) );
  AOI32V2_8TH40 U19 ( .A1(n97), .A2(n98), .A3(n99), .B1(B[6]), .B2(n13), .ZN(
        n96) );
  OAI21V2_8TH40 U20 ( .A1(A[5]), .A2(n29), .B(n100), .ZN(n99) );
  AOI32V2_8TH40 U21 ( .A1(n101), .A2(n69), .A3(n102), .B1(B[4]), .B2(n14), 
        .ZN(n100) );
  OAI21V2_8TH40 U22 ( .A1(A[17]), .A2(n23), .B(n85), .ZN(n84) );
  OAI21V2_8TH40 U23 ( .A1(A[11]), .A2(n26), .B(n91), .ZN(n90) );
  OAI21V2_8TH40 U24 ( .A1(A[23]), .A2(n20), .B(n79), .ZN(n78) );
  INV2_8TH40 U25 ( .I(A[1]), .ZN(n15) );
  INV2_8TH40 U26 ( .I(A[30]), .ZN(n1) );
  INV2_8TH40 U27 ( .I(A[10]), .ZN(n11) );
  INV2_8TH40 U28 ( .I(A[16]), .ZN(n8) );
  INV2_8TH40 U29 ( .I(A[22]), .ZN(n5) );
  INV2_8TH40 U30 ( .I(A[28]), .ZN(n2) );
  INV2_8TH40 U31 ( .I(A[18]), .ZN(n7) );
  INV2_8TH40 U32 ( .I(A[12]), .ZN(n10) );
  INV2_8TH40 U33 ( .I(A[24]), .ZN(n4) );
  INV2_8TH40 U34 ( .I(A[4]), .ZN(n14) );
  INV2_8TH40 U35 ( .I(A[14]), .ZN(n9) );
  INV2_8TH40 U36 ( .I(A[6]), .ZN(n13) );
  INV2_8TH40 U37 ( .I(A[8]), .ZN(n12) );
  INV2_8TH40 U38 ( .I(A[26]), .ZN(n3) );
  INV2_8TH40 U39 ( .I(B[31]), .ZN(n16) );
  INV2_8TH40 U40 ( .I(A[20]), .ZN(n6) );
  INV2_8TH40 U41 ( .I(B[17]), .ZN(n23) );
  INV2_8TH40 U42 ( .I(B[27]), .ZN(n18) );
  INV2_8TH40 U43 ( .I(B[29]), .ZN(n17) );
  INV2_8TH40 U44 ( .I(B[19]), .ZN(n22) );
  INV2_8TH40 U45 ( .I(B[5]), .ZN(n29) );
  INV2_8TH40 U46 ( .I(B[7]), .ZN(n28) );
  INV2_8TH40 U47 ( .I(B[9]), .ZN(n27) );
  INV2_8TH40 U48 ( .I(B[11]), .ZN(n26) );
  INV2_8TH40 U49 ( .I(B[23]), .ZN(n20) );
  INV2_8TH40 U50 ( .I(B[25]), .ZN(n19) );
  INV2_8TH40 U51 ( .I(B[15]), .ZN(n24) );
  INV2_8TH40 U52 ( .I(B[13]), .ZN(n25) );
  INV2_8TH40 U53 ( .I(B[3]), .ZN(n30) );
  INV2_8TH40 U54 ( .I(B[1]), .ZN(n32) );
  INV2_8TH40 U55 ( .I(B[2]), .ZN(n31) );
  INV2_8TH40 U56 ( .I(B[21]), .ZN(n21) );
  NAND4V0P5_8TH40 U57 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(n40) );
  OAI22V0_8TH40 U58 ( .A1(A[1]), .A2(n45), .B1(n45), .B2(n32), .ZN(n41) );
  INOR2V0_8TH40 U59 ( .A1(A[0]), .B1(B[0]), .ZN(n45) );
  NAND4V0P5_8TH40 U60 ( .A1(n46), .A2(n47), .A3(n48), .A4(n49), .ZN(n39) );
  NAND4V0P5_8TH40 U61 ( .A1(n50), .A2(n51), .A3(n52), .A4(n53), .ZN(n38) );
  NAND4V0P5_8TH40 U62 ( .A1(n54), .A2(n55), .A3(n56), .A4(n57), .ZN(n37) );
  NAND4V0P5_8TH40 U63 ( .A1(n60), .A2(n61), .A3(n62), .A4(n63), .ZN(n59) );
  NAND4V0P5_8TH40 U64 ( .A1(n64), .A2(n65), .A3(n66), .A4(n67), .ZN(n58) );
  I2NOR4V0_8TH40 U65 ( .A1(n68), .A2(n69), .B1(LT), .B2(n70), .ZN(n34) );
  OAI22V0_8TH40 U66 ( .A1(A[31]), .A2(n16), .B1(n70), .B2(n71), .ZN(LT) );
  AOI32V0_8TH40 U67 ( .A1(n44), .A2(n46), .A3(n74), .B1(B[28]), .B2(n2), .ZN(
        n73) );
  OAI21V0_8TH40 U68 ( .A1(A[25]), .A2(n19), .B(n77), .ZN(n76) );
  AOI32V0_8TH40 U69 ( .A1(n51), .A2(n52), .A3(n80), .B1(B[22]), .B2(n5), .ZN(
        n79) );
  OAI21V0_8TH40 U70 ( .A1(A[19]), .A2(n22), .B(n83), .ZN(n82) );
  AOI32V0_8TH40 U71 ( .A1(n57), .A2(n60), .A3(n86), .B1(B[16]), .B2(n8), .ZN(
        n85) );
  OAI21V0_8TH40 U72 ( .A1(A[13]), .A2(n25), .B(n89), .ZN(n88) );
  AOI32V0_8TH40 U73 ( .A1(n65), .A2(n66), .A3(n92), .B1(B[10]), .B2(n11), .ZN(
        n91) );
  OAI221V0_8TH40 U74 ( .A1(A[2]), .A2(n31), .B1(A[3]), .B2(n30), .C(n103), 
        .ZN(n102) );
  IOA21V0_8TH40 U75 ( .A1(n15), .A2(n104), .B(n32), .ZN(n105) );
  INOR2V0_8TH40 U76 ( .A1(B[0]), .B1(A[0]), .ZN(n104) );
  INAND2V0_8TH40 U77 ( .A1(B[8]), .B1(A[8]), .ZN(n67) );
  CLKNAND2V1_8TH40 U78 ( .A1(A[9]), .A2(n27), .ZN(n66) );
  INAND2V0_8TH40 U79 ( .A1(B[10]), .B1(A[10]), .ZN(n65) );
  CLKNAND2V1_8TH40 U80 ( .A1(A[11]), .A2(n26), .ZN(n64) );
  INAND2V0_8TH40 U81 ( .A1(B[12]), .B1(A[12]), .ZN(n63) );
  CLKNAND2V1_8TH40 U82 ( .A1(A[13]), .A2(n25), .ZN(n62) );
  INAND2V0_8TH40 U83 ( .A1(B[14]), .B1(A[14]), .ZN(n61) );
  CLKNAND2V1_8TH40 U84 ( .A1(A[15]), .A2(n24), .ZN(n60) );
  INAND2V0_8TH40 U85 ( .A1(B[16]), .B1(A[16]), .ZN(n57) );
  CLKNAND2V1_8TH40 U86 ( .A1(A[17]), .A2(n23), .ZN(n56) );
  INAND2V0_8TH40 U87 ( .A1(B[18]), .B1(A[18]), .ZN(n55) );
  CLKNAND2V1_8TH40 U88 ( .A1(A[19]), .A2(n22), .ZN(n54) );
  INAND2V0_8TH40 U89 ( .A1(B[20]), .B1(A[20]), .ZN(n53) );
  CLKNAND2V1_8TH40 U90 ( .A1(A[21]), .A2(n21), .ZN(n52) );
  INAND2V0_8TH40 U91 ( .A1(B[22]), .B1(A[22]), .ZN(n51) );
  CLKNAND2V1_8TH40 U92 ( .A1(A[23]), .A2(n20), .ZN(n50) );
  INAND2V0_8TH40 U93 ( .A1(B[24]), .B1(A[24]), .ZN(n49) );
  CLKNAND2V1_8TH40 U94 ( .A1(A[25]), .A2(n19), .ZN(n48) );
  INAND2V0_8TH40 U95 ( .A1(B[26]), .B1(A[26]), .ZN(n47) );
  CLKNAND2V1_8TH40 U96 ( .A1(A[27]), .A2(n18), .ZN(n46) );
  INAND2V0_8TH40 U97 ( .A1(B[28]), .B1(A[28]), .ZN(n44) );
  INAND2V0_8TH40 U98 ( .A1(B[30]), .B1(A[30]), .ZN(n43) );
  CLKNAND2V1_8TH40 U99 ( .A1(A[29]), .A2(n17), .ZN(n42) );
  AND2V0_8TH40 U100 ( .A1(A[31]), .A2(n16), .Z(n70) );
  CLKNAND2V1_8TH40 U101 ( .A1(A[3]), .A2(n30), .ZN(n69) );
  CLKNAND2V1_8TH40 U102 ( .A1(A[2]), .A2(n31), .ZN(n68) );
  AND4V0_8TH40 U103 ( .A1(n101), .A2(n98), .A3(n97), .A4(n94), .Z(n33) );
  CLKNAND2V1_8TH40 U104 ( .A1(A[7]), .A2(n28), .ZN(n94) );
  OR2V0_8TH40 U105 ( .A1(B[6]), .A2(n13), .Z(n97) );
  CLKNAND2V1_8TH40 U106 ( .A1(A[5]), .A2(n29), .ZN(n98) );
  OR2V0_8TH40 U107 ( .A1(B[4]), .A2(n14), .Z(n101) );
endmodule


module inst_execute ( rst, inst_type, inst_class, gpr1_data, gpr2_data, 
        target_gpr, gpr_we, hi_i, lo_i, df_wbex_hi, df_wbex_lo, 
        df_wbex_hilo_we, df_memex_hi, df_memex_lo, df_memex_hilo_we, 
        hilo_tmp_i, cycl_cnt_i, cur_inst_delayslot_i, link_addr, div_res, 
        div_done, inst_i, except_type_i, cur_inst_addr_i, hi_o, lo_o, hilo_we, 
        gpr_we_o, target_gpr_o, exe_result_o, hilo_tmp_o, cycl_cnt_o, 
        stall_req, signed_div, div_opdata1, div_opdata2, div_start, 
        inst_type_o, dmem_addr, ls_data_tmp, mem_cp0_we, mem_cp0_waddr, 
        mem_cp0_wdata, wb_cp0_we, wb_cp0_waddr, wb_cp0_wdata, cp0_ex_rdata, 
        ex_cp0_raddr, cp0_we, cp0_waddr, cp0_wdata, except_type_o, 
        cur_inst_addr_o, cur_inst_delayslot_o );
  input [7:0] inst_type;
  input [2:0] inst_class;
  input [31:0] gpr1_data;
  input [31:0] gpr2_data;
  input [4:0] target_gpr;
  input [31:0] hi_i;
  input [31:0] lo_i;
  input [31:0] df_wbex_hi;
  input [31:0] df_wbex_lo;
  input [31:0] df_memex_hi;
  input [31:0] df_memex_lo;
  input [63:0] hilo_tmp_i;
  input [1:0] cycl_cnt_i;
  input [31:0] link_addr;
  input [63:0] div_res;
  input [31:0] inst_i;
  input [31:0] except_type_i;
  input [31:0] cur_inst_addr_i;
  output [31:0] hi_o;
  output [31:0] lo_o;
  output [4:0] target_gpr_o;
  output [31:0] exe_result_o;
  output [63:0] hilo_tmp_o;
  output [1:0] cycl_cnt_o;
  output [31:0] div_opdata1;
  output [31:0] div_opdata2;
  output [7:0] inst_type_o;
  output [31:0] dmem_addr;
  output [31:0] ls_data_tmp;
  input [4:0] mem_cp0_waddr;
  input [31:0] mem_cp0_wdata;
  input [4:0] wb_cp0_waddr;
  input [31:0] wb_cp0_wdata;
  input [31:0] cp0_ex_rdata;
  output [4:0] ex_cp0_raddr;
  output [4:0] cp0_waddr;
  output [31:0] cp0_wdata;
  output [31:0] except_type_o;
  output [31:0] cur_inst_addr_o;
  input rst, gpr_we, df_wbex_hilo_we, df_memex_hilo_we, cur_inst_delayslot_i,
         div_done, mem_cp0_we, wb_cp0_we;
  output hilo_we, gpr_we_o, stall_req, signed_div, div_start, cp0_we,
         cur_inst_delayslot_o;
  wire   cur_inst_delayslot_i, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N96, N500, N501, N502,
         N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, N666, maddmsub_stall_req, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781,
         N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792,
         N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N818, N819, N951, N952, N953, N954, N955, N956,
         N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967,
         N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978,
         N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989,
         N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000,
         N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010,
         N1011, N1012, N1013, N1212, N1213, N1214, N1215, N1216, N1217, N1218,
         N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228,
         N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238,
         N1239, N1240, N1241, N1242, N1243, N1244, N1246, N1247, N1248, N1249,
         N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259,
         N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269,
         N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1348, N1349, N1350,
         N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360,
         N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370,
         N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380,
         N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390,
         N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400,
         N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410,
         N1411, N1412, N1413, N1414, N1416, N1574, N1807, N1808, N1809, N1810,
         N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820,
         N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1828, N1829, N1830,
         N1831, N1832, N1833, N1834, N1835, N1836, N1837, N1838, N1839, N1840,
         N1841, N1842, N1843, N1844, N1845, N1846, N1847, N1848, N1849, N1850,
         N1851, N1852, N1853, N1854, N1855, N1856, N1857, N1858, N1859, N1860,
         N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870,
         N1872, N1873, N1875, N2186, n1, n2, n3, n4, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         SYNOPSYS_UNCONNECTED_1;
  wire   [30:0] com_gpr2_data;
  wire   [31:0] sum_res;
  wire   [31:0] mul_opdata1;
  wire   [31:0] mul_opdata2;
  wire   [63:0] mul_res_tmp;
  wire   [31:0] lo;
  wire   [63:0] mul_res_tmp1;
  assign target_gpr_o[4] = target_gpr[4];
  assign target_gpr_o[3] = target_gpr[3];
  assign target_gpr_o[2] = target_gpr[2];
  assign target_gpr_o[1] = target_gpr[1];
  assign target_gpr_o[0] = target_gpr[0];
  assign inst_type_o[7] = inst_type[7];
  assign inst_type_o[6] = inst_type[6];
  assign inst_type_o[5] = inst_type[5];
  assign inst_type_o[4] = inst_type[4];
  assign inst_type_o[3] = inst_type[3];
  assign inst_type_o[2] = inst_type[2];
  assign inst_type_o[1] = inst_type[1];
  assign inst_type_o[0] = inst_type[0];
  assign ls_data_tmp[31] = gpr2_data[31];
  assign ls_data_tmp[30] = gpr2_data[30];
  assign ls_data_tmp[29] = gpr2_data[29];
  assign ls_data_tmp[28] = gpr2_data[28];
  assign ls_data_tmp[27] = gpr2_data[27];
  assign ls_data_tmp[26] = gpr2_data[26];
  assign ls_data_tmp[25] = gpr2_data[25];
  assign ls_data_tmp[24] = gpr2_data[24];
  assign ls_data_tmp[23] = gpr2_data[23];
  assign ls_data_tmp[22] = gpr2_data[22];
  assign ls_data_tmp[21] = gpr2_data[21];
  assign ls_data_tmp[20] = gpr2_data[20];
  assign ls_data_tmp[19] = gpr2_data[19];
  assign ls_data_tmp[18] = gpr2_data[18];
  assign ls_data_tmp[17] = gpr2_data[17];
  assign ls_data_tmp[16] = gpr2_data[16];
  assign ls_data_tmp[15] = gpr2_data[15];
  assign ls_data_tmp[14] = gpr2_data[14];
  assign ls_data_tmp[13] = gpr2_data[13];
  assign ls_data_tmp[12] = gpr2_data[12];
  assign ls_data_tmp[11] = gpr2_data[11];
  assign ls_data_tmp[10] = gpr2_data[10];
  assign ls_data_tmp[9] = gpr2_data[9];
  assign ls_data_tmp[8] = gpr2_data[8];
  assign ls_data_tmp[7] = gpr2_data[7];
  assign ls_data_tmp[6] = gpr2_data[6];
  assign ls_data_tmp[5] = gpr2_data[5];
  assign ls_data_tmp[4] = gpr2_data[4];
  assign ls_data_tmp[3] = gpr2_data[3];
  assign ls_data_tmp[2] = gpr2_data[2];
  assign ls_data_tmp[1] = gpr2_data[1];
  assign ls_data_tmp[0] = gpr2_data[0];
  assign except_type_o[12] = except_type_i[12];
  assign except_type_o[9] = except_type_i[9];
  assign except_type_o[8] = except_type_i[8];
  assign cur_inst_addr_o[31] = cur_inst_addr_i[31];
  assign cur_inst_addr_o[30] = cur_inst_addr_i[30];
  assign cur_inst_addr_o[29] = cur_inst_addr_i[29];
  assign cur_inst_addr_o[28] = cur_inst_addr_i[28];
  assign cur_inst_addr_o[27] = cur_inst_addr_i[27];
  assign cur_inst_addr_o[26] = cur_inst_addr_i[26];
  assign cur_inst_addr_o[25] = cur_inst_addr_i[25];
  assign cur_inst_addr_o[24] = cur_inst_addr_i[24];
  assign cur_inst_addr_o[23] = cur_inst_addr_i[23];
  assign cur_inst_addr_o[22] = cur_inst_addr_i[22];
  assign cur_inst_addr_o[21] = cur_inst_addr_i[21];
  assign cur_inst_addr_o[20] = cur_inst_addr_i[20];
  assign cur_inst_addr_o[19] = cur_inst_addr_i[19];
  assign cur_inst_addr_o[18] = cur_inst_addr_i[18];
  assign cur_inst_addr_o[17] = cur_inst_addr_i[17];
  assign cur_inst_addr_o[16] = cur_inst_addr_i[16];
  assign cur_inst_addr_o[15] = cur_inst_addr_i[15];
  assign cur_inst_addr_o[14] = cur_inst_addr_i[14];
  assign cur_inst_addr_o[13] = cur_inst_addr_i[13];
  assign cur_inst_addr_o[12] = cur_inst_addr_i[12];
  assign cur_inst_addr_o[11] = cur_inst_addr_i[11];
  assign cur_inst_addr_o[10] = cur_inst_addr_i[10];
  assign cur_inst_addr_o[9] = cur_inst_addr_i[9];
  assign cur_inst_addr_o[8] = cur_inst_addr_i[8];
  assign cur_inst_addr_o[7] = cur_inst_addr_i[7];
  assign cur_inst_addr_o[6] = cur_inst_addr_i[6];
  assign cur_inst_addr_o[5] = cur_inst_addr_i[5];
  assign cur_inst_addr_o[4] = cur_inst_addr_i[4];
  assign cur_inst_addr_o[3] = cur_inst_addr_i[3];
  assign cur_inst_addr_o[2] = cur_inst_addr_i[2];
  assign cur_inst_addr_o[1] = cur_inst_addr_i[1];
  assign cur_inst_addr_o[0] = cur_inst_addr_i[0];
  assign cur_inst_delayslot_o = cur_inst_delayslot_i;

  LAHQV1_8TH40 cycl_cnt_o_reg_1_ ( .E(N1413), .D(N1412), .Q(cycl_cnt_o[1]) );
  LAHQV1_8TH40 cycl_cnt_o_reg_0_ ( .E(N1413), .D(N1414), .Q(cycl_cnt_o[0]) );
  LAHQV1_8TH40 maddmsub_stall_req_reg ( .E(N1413), .D(N1414), .Q(
        maddmsub_stall_req) );
  LAHQV1_8TH40 ex_cp0_raddr_reg_4_ ( .E(N2186), .D(inst_i[15]), .Q(
        ex_cp0_raddr[4]) );
  LAHQV1_8TH40 ex_cp0_raddr_reg_3_ ( .E(N2186), .D(inst_i[14]), .Q(
        ex_cp0_raddr[3]) );
  LAHQV1_8TH40 ex_cp0_raddr_reg_2_ ( .E(N2186), .D(inst_i[13]), .Q(
        ex_cp0_raddr[2]) );
  LAHQV1_8TH40 ex_cp0_raddr_reg_1_ ( .E(N2186), .D(inst_i[12]), .Q(
        ex_cp0_raddr[1]) );
  LAHQV1_8TH40 ex_cp0_raddr_reg_0_ ( .E(N2186), .D(inst_i[11]), .Q(
        ex_cp0_raddr[0]) );
  inst_execute_DW01_ash_1 sll_482 ( .A(gpr2_data), .DATA_TC(1'b0), .SH(
        gpr1_data[4:0]), .SH_TC(1'b0), .B({N1838, N1837, N1836, N1835, N1834, 
        N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, 
        N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, 
        N1813, N1812, N1811, N1810, N1809, N1808, N1807}) );
  inst_execute_DW01_sub_1 sub_add_303_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
        n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
        n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
        n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
        n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
        n977, n978, n979, n980, n1013}), .CI(1'b0), .DIFF({N1013, N1012, N1011, 
        N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, 
        N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, 
        N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, 
        N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, 
        N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, 
        N953, N952, N951, SYNOPSYS_UNCONNECTED_1}) );
  inst_execute_DW01_sub_2 sub_add_260_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B(mul_res_tmp), .CI(1'b0), .DIFF({N666, N665, N664, N663, N662, N661, 
        N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, 
        N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, 
        N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, 
        N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, 
        N612, N611, N610, N609, N608, N607, N606, N605, N604, N603}) );
  inst_execute_DW02_mult_0 mult_243 ( .A(mul_opdata1), .B(mul_opdata2), .TC(
        1'b0), .PRODUCT(mul_res_tmp) );
  inst_execute_DW01_inc_0 add_237 ( .A({n1042, n1043, n1044, n1045, n1046, 
        n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
        n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
        n1067, n1068, n1069, n1070, n1071, n1072, n1073}), .SUM({N596, N595, 
        N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, 
        N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, 
        N570, N569, N568, N567, N566, N565}) );
  inst_execute_DW01_inc_1 add_230 ( .A({n1015, n1016, n1017, n1018, n1019, 
        n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
        n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
        n1040, n1041, n916, n915, n914, n913, n912}), .SUM({N531, N530, N529, 
        N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, 
        N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, 
        N504, N503, N502, N501, N500}) );
  inst_execute_DW01_add_1 add_139 ( .A(gpr1_data), .B({n917, com_gpr2_data}), 
        .CI(1'b0), .SUM(sum_res) );
  inst_execute_DW01_sub_3 sub_add_127_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(gpr2_data), .CI(1'b0), .DIFF({N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, 
        N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, 
        N60}) );
  inst_execute_DW01_add_2 add_118 ( .A(gpr1_data), .B({inst_i[15], inst_i[15], 
        inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], 
        inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], inst_i[15], 
        inst_i[15], inst_i[15], inst_i[15:0]}), .CI(1'b0), .SUM(dmem_addr) );
  inst_execute_DW_rash_0 r204 ( .A(gpr2_data), .DATA_TC(1'b0), .SH(
        gpr1_data[4:0]), .SH_TC(1'b0), .B({N1870, N1869, N1868, N1867, N1866, 
        N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, 
        N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, 
        N1845, N1844, N1843, N1842, N1841, N1840, N1839}) );
  inst_execute_DW01_add_3 r201 ( .A(hilo_tmp_i), .B({n981, n982, n983, n984, 
        n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
        n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
        n1007, n1008, n1009, n1010, n1011, n1012, lo}), .CI(1'b0), .SUM({N819, 
        N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, 
        N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, 
        N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, 
        N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, 
        N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, 
        N758, N757, N756}) );
  inst_execute_DW01_cmp6_2 r196 ( .A(gpr1_data), .B(gpr2_data), .TC(1'b0), 
        .LT(N96), .NE(N1574) );
  LAHQV4_8TH40 mul_res_tmp1_reg_63_ ( .E(N1416), .D(N1276), .Q(
        mul_res_tmp1[63]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_62_ ( .E(N1416), .D(N1275), .Q(
        mul_res_tmp1[62]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_61_ ( .E(N1416), .D(N1274), .Q(
        mul_res_tmp1[61]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_60_ ( .E(N1416), .D(N1273), .Q(
        mul_res_tmp1[60]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_59_ ( .E(N1416), .D(N1272), .Q(
        mul_res_tmp1[59]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_58_ ( .E(N1416), .D(N1271), .Q(
        mul_res_tmp1[58]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_57_ ( .E(N1416), .D(N1270), .Q(
        mul_res_tmp1[57]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_56_ ( .E(N1416), .D(N1269), .Q(
        mul_res_tmp1[56]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_55_ ( .E(N1416), .D(N1268), .Q(
        mul_res_tmp1[55]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_54_ ( .E(N1416), .D(N1267), .Q(
        mul_res_tmp1[54]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_53_ ( .E(N1416), .D(N1266), .Q(
        mul_res_tmp1[53]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_52_ ( .E(N1416), .D(N1265), .Q(
        mul_res_tmp1[52]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_51_ ( .E(N1416), .D(N1264), .Q(
        mul_res_tmp1[51]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_50_ ( .E(N1416), .D(N1263), .Q(
        mul_res_tmp1[50]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_49_ ( .E(N1416), .D(N1262), .Q(
        mul_res_tmp1[49]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_48_ ( .E(N1416), .D(N1261), .Q(
        mul_res_tmp1[48]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_47_ ( .E(N1416), .D(N1260), .Q(
        mul_res_tmp1[47]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_46_ ( .E(N1416), .D(N1259), .Q(
        mul_res_tmp1[46]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_45_ ( .E(N1416), .D(N1258), .Q(
        mul_res_tmp1[45]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_44_ ( .E(N1416), .D(N1257), .Q(
        mul_res_tmp1[44]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_43_ ( .E(N1416), .D(N1256), .Q(
        mul_res_tmp1[43]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_42_ ( .E(N1416), .D(N1255), .Q(
        mul_res_tmp1[42]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_41_ ( .E(N1416), .D(N1254), .Q(
        mul_res_tmp1[41]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_40_ ( .E(N1416), .D(N1253), .Q(
        mul_res_tmp1[40]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_39_ ( .E(N1416), .D(N1252), .Q(
        mul_res_tmp1[39]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_38_ ( .E(N1416), .D(N1251), .Q(
        mul_res_tmp1[38]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_37_ ( .E(N1416), .D(N1250), .Q(
        mul_res_tmp1[37]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_36_ ( .E(N1416), .D(N1249), .Q(
        mul_res_tmp1[36]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_35_ ( .E(N1416), .D(N1248), .Q(
        mul_res_tmp1[35]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_34_ ( .E(N1416), .D(N1247), .Q(
        mul_res_tmp1[34]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_33_ ( .E(N1416), .D(N1246), .Q(
        mul_res_tmp1[33]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_32_ ( .E(N1416), .D(N1244), .Q(
        mul_res_tmp1[32]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_31_ ( .E(N1416), .D(N1243), .Q(
        mul_res_tmp1[31]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_30_ ( .E(N1416), .D(N1242), .Q(
        mul_res_tmp1[30]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_29_ ( .E(N1416), .D(N1241), .Q(
        mul_res_tmp1[29]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_28_ ( .E(N1416), .D(N1240), .Q(
        mul_res_tmp1[28]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_27_ ( .E(N1416), .D(N1239), .Q(
        mul_res_tmp1[27]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_26_ ( .E(N1416), .D(N1238), .Q(
        mul_res_tmp1[26]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_25_ ( .E(N1416), .D(N1237), .Q(
        mul_res_tmp1[25]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_24_ ( .E(N1416), .D(N1236), .Q(
        mul_res_tmp1[24]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_23_ ( .E(N1416), .D(N1235), .Q(
        mul_res_tmp1[23]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_22_ ( .E(N1416), .D(N1234), .Q(
        mul_res_tmp1[22]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_21_ ( .E(N1416), .D(N1233), .Q(
        mul_res_tmp1[21]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_20_ ( .E(N1416), .D(N1232), .Q(
        mul_res_tmp1[20]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_19_ ( .E(N1416), .D(N1231), .Q(
        mul_res_tmp1[19]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_18_ ( .E(N1416), .D(N1230), .Q(
        mul_res_tmp1[18]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_17_ ( .E(N1416), .D(N1229), .Q(
        mul_res_tmp1[17]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_16_ ( .E(N1416), .D(N1228), .Q(
        mul_res_tmp1[16]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_15_ ( .E(N1416), .D(N1227), .Q(
        mul_res_tmp1[15]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_14_ ( .E(N1416), .D(N1226), .Q(
        mul_res_tmp1[14]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_13_ ( .E(N1416), .D(N1225), .Q(
        mul_res_tmp1[13]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_12_ ( .E(N1416), .D(N1224), .Q(
        mul_res_tmp1[12]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_11_ ( .E(N1416), .D(N1223), .Q(
        mul_res_tmp1[11]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_10_ ( .E(N1416), .D(N1222), .Q(
        mul_res_tmp1[10]) );
  LAHQV4_8TH40 mul_res_tmp1_reg_9_ ( .E(N1416), .D(N1221), .Q(mul_res_tmp1[9])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_8_ ( .E(N1416), .D(N1220), .Q(mul_res_tmp1[8])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_7_ ( .E(N1416), .D(N1219), .Q(mul_res_tmp1[7])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_6_ ( .E(N1416), .D(N1218), .Q(mul_res_tmp1[6])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_5_ ( .E(N1416), .D(N1217), .Q(mul_res_tmp1[5])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_4_ ( .E(N1416), .D(N1216), .Q(mul_res_tmp1[4])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_3_ ( .E(N1416), .D(N1215), .Q(mul_res_tmp1[3])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_2_ ( .E(N1416), .D(N1214), .Q(mul_res_tmp1[2])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_1_ ( .E(N1416), .D(N1213), .Q(mul_res_tmp1[1])
         );
  LAHQV4_8TH40 mul_res_tmp1_reg_0_ ( .E(N1416), .D(N1212), .Q(mul_res_tmp1[0])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_63_ ( .E(N1413), .D(N1411), .Q(hilo_tmp_o[63])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_62_ ( .E(N1413), .D(N1410), .Q(hilo_tmp_o[62])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_61_ ( .E(N1413), .D(N1409), .Q(hilo_tmp_o[61])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_60_ ( .E(N1413), .D(N1408), .Q(hilo_tmp_o[60])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_59_ ( .E(N1413), .D(N1407), .Q(hilo_tmp_o[59])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_58_ ( .E(N1413), .D(N1406), .Q(hilo_tmp_o[58])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_57_ ( .E(N1413), .D(N1405), .Q(hilo_tmp_o[57])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_56_ ( .E(N1413), .D(N1404), .Q(hilo_tmp_o[56])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_55_ ( .E(N1413), .D(N1403), .Q(hilo_tmp_o[55])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_54_ ( .E(N1413), .D(N1402), .Q(hilo_tmp_o[54])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_53_ ( .E(N1413), .D(N1401), .Q(hilo_tmp_o[53])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_52_ ( .E(N1413), .D(N1400), .Q(hilo_tmp_o[52])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_51_ ( .E(N1413), .D(N1399), .Q(hilo_tmp_o[51])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_50_ ( .E(N1413), .D(N1398), .Q(hilo_tmp_o[50])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_49_ ( .E(N1413), .D(N1397), .Q(hilo_tmp_o[49])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_48_ ( .E(N1413), .D(N1396), .Q(hilo_tmp_o[48])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_47_ ( .E(N1413), .D(N1395), .Q(hilo_tmp_o[47])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_46_ ( .E(N1413), .D(N1394), .Q(hilo_tmp_o[46])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_45_ ( .E(N1413), .D(N1393), .Q(hilo_tmp_o[45])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_44_ ( .E(N1413), .D(N1392), .Q(hilo_tmp_o[44])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_43_ ( .E(N1413), .D(N1391), .Q(hilo_tmp_o[43])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_42_ ( .E(N1413), .D(N1390), .Q(hilo_tmp_o[42])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_41_ ( .E(N1413), .D(N1389), .Q(hilo_tmp_o[41])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_40_ ( .E(N1413), .D(N1388), .Q(hilo_tmp_o[40])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_39_ ( .E(N1413), .D(N1387), .Q(hilo_tmp_o[39])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_38_ ( .E(N1413), .D(N1386), .Q(hilo_tmp_o[38])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_37_ ( .E(N1413), .D(N1385), .Q(hilo_tmp_o[37])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_36_ ( .E(N1413), .D(N1384), .Q(hilo_tmp_o[36])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_35_ ( .E(N1413), .D(N1383), .Q(hilo_tmp_o[35])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_34_ ( .E(N1413), .D(N1382), .Q(hilo_tmp_o[34])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_33_ ( .E(N1413), .D(N1381), .Q(hilo_tmp_o[33])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_32_ ( .E(N1413), .D(N1380), .Q(hilo_tmp_o[32])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_31_ ( .E(N1413), .D(N1379), .Q(hilo_tmp_o[31])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_30_ ( .E(N1413), .D(N1378), .Q(hilo_tmp_o[30])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_29_ ( .E(N1413), .D(N1377), .Q(hilo_tmp_o[29])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_28_ ( .E(N1413), .D(N1376), .Q(hilo_tmp_o[28])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_27_ ( .E(N1413), .D(N1375), .Q(hilo_tmp_o[27])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_26_ ( .E(N1413), .D(N1374), .Q(hilo_tmp_o[26])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_25_ ( .E(N1413), .D(N1373), .Q(hilo_tmp_o[25])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_24_ ( .E(N1413), .D(N1372), .Q(hilo_tmp_o[24])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_23_ ( .E(N1413), .D(N1371), .Q(hilo_tmp_o[23])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_22_ ( .E(N1413), .D(N1370), .Q(hilo_tmp_o[22])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_21_ ( .E(N1413), .D(N1369), .Q(hilo_tmp_o[21])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_20_ ( .E(N1413), .D(N1368), .Q(hilo_tmp_o[20])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_19_ ( .E(N1413), .D(N1367), .Q(hilo_tmp_o[19])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_18_ ( .E(N1413), .D(N1366), .Q(hilo_tmp_o[18])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_17_ ( .E(N1413), .D(N1365), .Q(hilo_tmp_o[17])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_16_ ( .E(N1413), .D(N1364), .Q(hilo_tmp_o[16])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_15_ ( .E(N1413), .D(N1363), .Q(hilo_tmp_o[15])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_14_ ( .E(N1413), .D(N1362), .Q(hilo_tmp_o[14])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_13_ ( .E(N1413), .D(N1361), .Q(hilo_tmp_o[13])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_12_ ( .E(N1413), .D(N1360), .Q(hilo_tmp_o[12])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_11_ ( .E(N1413), .D(N1359), .Q(hilo_tmp_o[11])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_10_ ( .E(N1413), .D(N1358), .Q(hilo_tmp_o[10])
         );
  LAHQV4_8TH40 hilo_tmp_o_reg_9_ ( .E(N1413), .D(N1357), .Q(hilo_tmp_o[9]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_8_ ( .E(N1413), .D(N1356), .Q(hilo_tmp_o[8]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_7_ ( .E(N1413), .D(N1355), .Q(hilo_tmp_o[7]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_6_ ( .E(N1413), .D(N1354), .Q(hilo_tmp_o[6]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_5_ ( .E(N1413), .D(N1353), .Q(hilo_tmp_o[5]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_4_ ( .E(N1413), .D(N1352), .Q(hilo_tmp_o[4]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_3_ ( .E(N1413), .D(N1351), .Q(hilo_tmp_o[3]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_2_ ( .E(N1413), .D(N1350), .Q(hilo_tmp_o[2]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_1_ ( .E(N1413), .D(N1349), .Q(hilo_tmp_o[1]) );
  LAHQV4_8TH40 hilo_tmp_o_reg_0_ ( .E(N1413), .D(N1348), .Q(hilo_tmp_o[0]) );
  AO211V2_8TH40 U3 ( .A1(n794), .A2(n839), .B(rst), .C(n840), .Z(n1) );
  XNOR2V2_8TH40 U4 ( .A1(n15), .A2(n915), .ZN(n2) );
  I2NAND4V2_8TH40 U5 ( .A1(cycl_cnt_i[0]), .A2(n840), .B1(n910), .B2(n777), 
        .ZN(n838) );
  NAND4V2_8TH40 U6 ( .A1(inst_type[0]), .A2(n234), .A3(n235), .A4(inst_type[1]), .ZN(n37) );
  INV2_8TH40 U7 ( .I(n1), .ZN(n3) );
  AOI21V4_8TH40 U8 ( .A1(n910), .A2(cycl_cnt_i[0]), .B(n759), .ZN(n911) );
  INOR2V4_8TH40 U9 ( .A1(N758), .B1(n911), .ZN(N1214) );
  INOR2V4_8TH40 U10 ( .A1(N759), .B1(n911), .ZN(N1215) );
  INOR2V4_8TH40 U11 ( .A1(N760), .B1(n911), .ZN(N1216) );
  INOR2V4_8TH40 U12 ( .A1(N761), .B1(n911), .ZN(N1217) );
  INOR2V4_8TH40 U13 ( .A1(N762), .B1(n911), .ZN(N1218) );
  INOR2V4_8TH40 U14 ( .A1(N763), .B1(n911), .ZN(N1219) );
  INOR2V4_8TH40 U15 ( .A1(N764), .B1(n911), .ZN(N1220) );
  INOR2V4_8TH40 U16 ( .A1(N765), .B1(n911), .ZN(N1221) );
  INOR2V4_8TH40 U17 ( .A1(N766), .B1(n911), .ZN(N1222) );
  INOR2V4_8TH40 U18 ( .A1(N767), .B1(n911), .ZN(N1223) );
  INOR2V4_8TH40 U19 ( .A1(N768), .B1(n911), .ZN(N1224) );
  INOR2V4_8TH40 U20 ( .A1(N769), .B1(n911), .ZN(N1225) );
  INOR2V4_8TH40 U21 ( .A1(N770), .B1(n911), .ZN(N1226) );
  INOR2V4_8TH40 U32 ( .A1(N771), .B1(n911), .ZN(N1227) );
  INOR2V4_8TH40 U33 ( .A1(N772), .B1(n911), .ZN(N1228) );
  INOR2V4_8TH40 U34 ( .A1(N773), .B1(n911), .ZN(N1229) );
  INOR2V4_8TH40 U35 ( .A1(N774), .B1(n911), .ZN(N1230) );
  INOR2V4_8TH40 U36 ( .A1(N775), .B1(n911), .ZN(N1231) );
  INOR2V4_8TH40 U37 ( .A1(N776), .B1(n911), .ZN(N1232) );
  INOR2V4_8TH40 U38 ( .A1(N777), .B1(n911), .ZN(N1233) );
  INOR2V4_8TH40 U39 ( .A1(N778), .B1(n911), .ZN(N1234) );
  INOR2V4_8TH40 U40 ( .A1(N779), .B1(n911), .ZN(N1235) );
  INOR2V4_8TH40 U41 ( .A1(N780), .B1(n911), .ZN(N1236) );
  INOR2V4_8TH40 U42 ( .A1(N781), .B1(n911), .ZN(N1237) );
  INOR2V4_8TH40 U43 ( .A1(N782), .B1(n911), .ZN(N1238) );
  INOR2V4_8TH40 U44 ( .A1(N783), .B1(n911), .ZN(N1239) );
  INOR2V4_8TH40 U45 ( .A1(N784), .B1(n911), .ZN(N1240) );
  INOR2V4_8TH40 U46 ( .A1(N785), .B1(n911), .ZN(N1241) );
  INOR2V4_8TH40 U47 ( .A1(N786), .B1(n911), .ZN(N1242) );
  INOR2V4_8TH40 U48 ( .A1(N787), .B1(n911), .ZN(N1243) );
  INOR2V4_8TH40 U49 ( .A1(N788), .B1(n911), .ZN(N1244) );
  INOR2V4_8TH40 U50 ( .A1(N789), .B1(n911), .ZN(N1246) );
  INOR2V4_8TH40 U51 ( .A1(N790), .B1(n911), .ZN(N1247) );
  INOR2V4_8TH40 U52 ( .A1(N791), .B1(n911), .ZN(N1248) );
  INOR2V4_8TH40 U53 ( .A1(N792), .B1(n911), .ZN(N1249) );
  INOR2V4_8TH40 U54 ( .A1(N793), .B1(n911), .ZN(N1250) );
  INOR2V4_8TH40 U55 ( .A1(N794), .B1(n911), .ZN(N1251) );
  INOR2V4_8TH40 U56 ( .A1(N795), .B1(n911), .ZN(N1252) );
  INOR2V4_8TH40 U57 ( .A1(N796), .B1(n911), .ZN(N1253) );
  INOR2V4_8TH40 U58 ( .A1(N797), .B1(n911), .ZN(N1254) );
  INOR2V4_8TH40 U59 ( .A1(N798), .B1(n911), .ZN(N1255) );
  INOR2V4_8TH40 U60 ( .A1(N799), .B1(n911), .ZN(N1256) );
  INOR2V4_8TH40 U61 ( .A1(N800), .B1(n911), .ZN(N1257) );
  INOR2V4_8TH40 U62 ( .A1(N801), .B1(n911), .ZN(N1258) );
  INOR2V4_8TH40 U63 ( .A1(N802), .B1(n911), .ZN(N1259) );
  INOR2V4_8TH40 U64 ( .A1(N803), .B1(n911), .ZN(N1260) );
  INOR2V4_8TH40 U65 ( .A1(N804), .B1(n911), .ZN(N1261) );
  INOR2V4_8TH40 U66 ( .A1(N805), .B1(n911), .ZN(N1262) );
  INOR2V4_8TH40 U67 ( .A1(N806), .B1(n911), .ZN(N1263) );
  INOR2V4_8TH40 U68 ( .A1(N807), .B1(n911), .ZN(N1264) );
  INOR2V4_8TH40 U69 ( .A1(N808), .B1(n911), .ZN(N1265) );
  INOR2V4_8TH40 U70 ( .A1(N809), .B1(n911), .ZN(N1266) );
  INOR2V4_8TH40 U71 ( .A1(N810), .B1(n911), .ZN(N1267) );
  INOR2V4_8TH40 U72 ( .A1(N811), .B1(n911), .ZN(N1268) );
  INOR2V4_8TH40 U73 ( .A1(N812), .B1(n911), .ZN(N1269) );
  INOR2V4_8TH40 U74 ( .A1(N813), .B1(n911), .ZN(N1270) );
  INOR2V4_8TH40 U75 ( .A1(N814), .B1(n911), .ZN(N1271) );
  INOR2V4_8TH40 U76 ( .A1(N815), .B1(n911), .ZN(N1272) );
  INOR2V4_8TH40 U77 ( .A1(N816), .B1(n911), .ZN(N1273) );
  INOR2V4_8TH40 U78 ( .A1(N817), .B1(n911), .ZN(N1274) );
  INOR2V4_8TH40 U79 ( .A1(N818), .B1(n911), .ZN(N1275) );
  INOR2V4_8TH40 U80 ( .A1(N819), .B1(n911), .ZN(N1276) );
  INOR2V4_8TH40 U81 ( .A1(N757), .B1(n911), .ZN(N1213) );
  INOR2V4_8TH40 U82 ( .A1(N756), .B1(n911), .ZN(N1212) );
  AOI22V2_8TH40 U83 ( .A1(n289), .A2(n983), .B1(cp0_ex_rdata[29]), .B2(n254), 
        .ZN(n474) );
  AOI22V2_8TH40 U84 ( .A1(n289), .A2(n985), .B1(cp0_ex_rdata[27]), .B2(n254), 
        .ZN(n498) );
  AOI22V2_8TH40 U85 ( .A1(n289), .A2(n986), .B1(cp0_ex_rdata[26]), .B2(n254), 
        .ZN(n510) );
  AOI22V2_8TH40 U86 ( .A1(n289), .A2(n987), .B1(cp0_ex_rdata[25]), .B2(n254), 
        .ZN(n521) );
  AOI22V2_8TH40 U87 ( .A1(n289), .A2(n988), .B1(cp0_ex_rdata[24]), .B2(n254), 
        .ZN(n533) );
  AOI22V2_8TH40 U88 ( .A1(n289), .A2(n990), .B1(cp0_ex_rdata[22]), .B2(n254), 
        .ZN(n556) );
  AOI22V2_8TH40 U89 ( .A1(n289), .A2(n992), .B1(cp0_ex_rdata[20]), .B2(n254), 
        .ZN(n578) );
  OAI22V2_8TH40 U90 ( .A1(n568), .A2(n838), .B1(n886), .B2(n842), .ZN(N1369)
         );
  OAI22V2_8TH40 U91 ( .A1(n149), .A2(n838), .B1(n841), .B2(n842), .ZN(N1411)
         );
  OAI22V2_8TH40 U92 ( .A1(n584), .A2(n838), .B1(n887), .B2(n842), .ZN(N1368)
         );
  OAI22V2_8TH40 U93 ( .A1(n633), .A2(n838), .B1(n888), .B2(n842), .ZN(N1367)
         );
  OAI22V2_8TH40 U94 ( .A1(n644), .A2(n838), .B1(n889), .B2(n842), .ZN(N1366)
         );
  OAI22V2_8TH40 U95 ( .A1(n654), .A2(n838), .B1(n890), .B2(n842), .ZN(N1365)
         );
  OAI22V2_8TH40 U96 ( .A1(n665), .A2(n838), .B1(n891), .B2(n842), .ZN(N1364)
         );
  OAI22V2_8TH40 U97 ( .A1(n675), .A2(n838), .B1(n892), .B2(n842), .ZN(N1363)
         );
  OAI22V2_8TH40 U98 ( .A1(n690), .A2(n838), .B1(n893), .B2(n842), .ZN(N1362)
         );
  OAI22V2_8TH40 U99 ( .A1(n697), .A2(n838), .B1(n894), .B2(n842), .ZN(N1361)
         );
  OAI22V2_8TH40 U100 ( .A1(n711), .A2(n838), .B1(n895), .B2(n842), .ZN(N1360)
         );
  OAI22V2_8TH40 U101 ( .A1(n717), .A2(n838), .B1(n896), .B2(n842), .ZN(N1359)
         );
  OAI22V2_8TH40 U102 ( .A1(n728), .A2(n838), .B1(n897), .B2(n842), .ZN(N1358)
         );
  OAI22V2_8TH40 U103 ( .A1(n253), .A2(n838), .B1(n898), .B2(n842), .ZN(N1357)
         );
  OAI22V2_8TH40 U104 ( .A1(n277), .A2(n838), .B1(n899), .B2(n842), .ZN(N1356)
         );
  OAI22V2_8TH40 U105 ( .A1(n287), .A2(n838), .B1(n900), .B2(n842), .ZN(N1355)
         );
  OAI22V2_8TH40 U106 ( .A1(n301), .A2(n838), .B1(n901), .B2(n842), .ZN(N1354)
         );
  OAI22V2_8TH40 U107 ( .A1(n330), .A2(n838), .B1(n902), .B2(n842), .ZN(N1353)
         );
  OAI22V2_8TH40 U108 ( .A1(n362), .A2(n838), .B1(n903), .B2(n842), .ZN(N1352)
         );
  OAI22V2_8TH40 U109 ( .A1(n391), .A2(n838), .B1(n904), .B2(n842), .ZN(N1351)
         );
  OAI22V2_8TH40 U110 ( .A1(n468), .A2(n838), .B1(n905), .B2(n842), .ZN(N1350)
         );
  OAI22V2_8TH40 U111 ( .A1(n627), .A2(n838), .B1(n906), .B2(n842), .ZN(N1349)
         );
  AOI22V2_8TH40 U112 ( .A1(n289), .A2(n1007), .B1(cp0_ex_rdata[5]), .B2(n254), 
        .ZN(n311) );
  MUX2NV2_8TH40 U113 ( .I0(n832), .I1(n833), .S(gpr1_data[31]), .ZN(n828) );
  AOI22V2_8TH40 U114 ( .A1(N1838), .A2(n262), .B1(n415), .B2(gpr2_data[31]), 
        .ZN(n410) );
  AOI22V2_8TH40 U115 ( .A1(wb_cp0_wdata[29]), .A2(n255), .B1(N1836), .B2(n262), 
        .ZN(n473) );
  AOI22V2_8TH40 U116 ( .A1(wb_cp0_wdata[27]), .A2(n255), .B1(N1834), .B2(n262), 
        .ZN(n497) );
  AOI22V2_8TH40 U117 ( .A1(wb_cp0_wdata[26]), .A2(n255), .B1(N1833), .B2(n262), 
        .ZN(n509) );
  AOI22V2_8TH40 U118 ( .A1(wb_cp0_wdata[25]), .A2(n255), .B1(N1832), .B2(n262), 
        .ZN(n520) );
  AOI22V2_8TH40 U119 ( .A1(wb_cp0_wdata[24]), .A2(n255), .B1(N1831), .B2(n262), 
        .ZN(n532) );
  AOI22V2_8TH40 U120 ( .A1(wb_cp0_wdata[22]), .A2(n255), .B1(N1829), .B2(n262), 
        .ZN(n555) );
  AOI22V2_8TH40 U121 ( .A1(wb_cp0_wdata[20]), .A2(n255), .B1(N1827), .B2(n262), 
        .ZN(n577) );
  AOI22V2_8TH40 U122 ( .A1(N1821), .A2(n262), .B1(n263), .B2(gpr1_data[14]), 
        .ZN(n683) );
  AOI22V2_8TH40 U123 ( .A1(N1819), .A2(n262), .B1(n263), .B2(gpr1_data[12]), 
        .ZN(n706) );
  OAI211V2_8TH40 U124 ( .A1(n1037), .A2(n37), .B(n38), .C(n39), .ZN(lo_o[9])
         );
  OAI211V2_8TH40 U125 ( .A1(n1038), .A2(n37), .B(n43), .C(n44), .ZN(lo_o[8])
         );
  OAI211V2_8TH40 U126 ( .A1(n1039), .A2(n37), .B(n45), .C(n46), .ZN(lo_o[7])
         );
  OAI211V2_8TH40 U127 ( .A1(n1040), .A2(n37), .B(n47), .C(n48), .ZN(lo_o[6])
         );
  OAI211V2_8TH40 U128 ( .A1(n1041), .A2(n37), .B(n49), .C(n50), .ZN(lo_o[5])
         );
  OAI211V2_8TH40 U129 ( .A1(n916), .A2(n37), .B(n51), .C(n52), .ZN(lo_o[4]) );
  OAI211V2_8TH40 U130 ( .A1(n915), .A2(n37), .B(n53), .C(n54), .ZN(lo_o[3]) );
  OAI211V2_8TH40 U131 ( .A1(n1015), .A2(n37), .B(n55), .C(n56), .ZN(lo_o[31])
         );
  OAI211V2_8TH40 U132 ( .A1(n1016), .A2(n37), .B(n57), .C(n58), .ZN(lo_o[30])
         );
  OAI211V2_8TH40 U133 ( .A1(n914), .A2(n37), .B(n59), .C(n60), .ZN(lo_o[2]) );
  OAI211V2_8TH40 U134 ( .A1(n1017), .A2(n37), .B(n61), .C(n62), .ZN(lo_o[29])
         );
  OAI211V2_8TH40 U135 ( .A1(n1018), .A2(n37), .B(n63), .C(n64), .ZN(lo_o[28])
         );
  OAI211V2_8TH40 U136 ( .A1(n1019), .A2(n37), .B(n65), .C(n66), .ZN(lo_o[27])
         );
  OAI211V2_8TH40 U137 ( .A1(n1020), .A2(n37), .B(n67), .C(n68), .ZN(lo_o[26])
         );
  OAI211V2_8TH40 U138 ( .A1(n1021), .A2(n37), .B(n69), .C(n70), .ZN(lo_o[25])
         );
  OAI211V2_8TH40 U139 ( .A1(n1022), .A2(n37), .B(n71), .C(n72), .ZN(lo_o[24])
         );
  OAI211V2_8TH40 U140 ( .A1(n1023), .A2(n37), .B(n73), .C(n74), .ZN(lo_o[23])
         );
  OAI211V2_8TH40 U141 ( .A1(n1024), .A2(n37), .B(n75), .C(n76), .ZN(lo_o[22])
         );
  OAI211V2_8TH40 U142 ( .A1(n1025), .A2(n37), .B(n77), .C(n78), .ZN(lo_o[21])
         );
  OAI211V2_8TH40 U143 ( .A1(n1026), .A2(n37), .B(n79), .C(n80), .ZN(lo_o[20])
         );
  OAI211V2_8TH40 U144 ( .A1(n913), .A2(n37), .B(n81), .C(n82), .ZN(lo_o[1]) );
  OAI211V2_8TH40 U145 ( .A1(n1027), .A2(n37), .B(n83), .C(n84), .ZN(lo_o[19])
         );
  OAI211V2_8TH40 U146 ( .A1(n1028), .A2(n37), .B(n85), .C(n86), .ZN(lo_o[18])
         );
  OAI211V2_8TH40 U147 ( .A1(n1029), .A2(n37), .B(n87), .C(n88), .ZN(lo_o[17])
         );
  OAI211V2_8TH40 U148 ( .A1(n1030), .A2(n37), .B(n89), .C(n90), .ZN(lo_o[16])
         );
  OAI211V2_8TH40 U149 ( .A1(n1031), .A2(n37), .B(n91), .C(n92), .ZN(lo_o[15])
         );
  OAI211V2_8TH40 U150 ( .A1(n1032), .A2(n37), .B(n93), .C(n94), .ZN(lo_o[14])
         );
  OAI211V2_8TH40 U151 ( .A1(n1033), .A2(n37), .B(n95), .C(n96), .ZN(lo_o[13])
         );
  OAI211V2_8TH40 U152 ( .A1(n1034), .A2(n37), .B(n97), .C(n98), .ZN(lo_o[12])
         );
  OAI211V2_8TH40 U153 ( .A1(n1035), .A2(n37), .B(n99), .C(n100), .ZN(lo_o[11])
         );
  OAI211V2_8TH40 U154 ( .A1(n1036), .A2(n37), .B(n101), .C(n102), .ZN(lo_o[10]) );
  OAI211V2_8TH40 U155 ( .A1(n912), .A2(n37), .B(n103), .C(n104), .ZN(lo_o[0])
         );
  NAND4V2S_8TH40 U156 ( .A1(n120), .A2(n37), .A3(n121), .A4(n18), .ZN(hilo_we)
         );
  OAI211V2_8TH40 U157 ( .A1(n28), .A2(n37), .B(n122), .C(n123), .ZN(hi_o[9])
         );
  OAI211V2_8TH40 U158 ( .A1(n29), .A2(n37), .B(n125), .C(n126), .ZN(hi_o[8])
         );
  OAI211V2_8TH40 U159 ( .A1(n128), .A2(n37), .B(n129), .C(n130), .ZN(hi_o[7])
         );
  OAI211V2_8TH40 U160 ( .A1(n30), .A2(n37), .B(n132), .C(n133), .ZN(hi_o[6])
         );
  OAI211V2_8TH40 U161 ( .A1(n135), .A2(n37), .B(n136), .C(n137), .ZN(hi_o[5])
         );
  OAI211V2_8TH40 U162 ( .A1(n31), .A2(n37), .B(n139), .C(n140), .ZN(hi_o[4])
         );
  OAI211V2_8TH40 U163 ( .A1(n142), .A2(n37), .B(n143), .C(n144), .ZN(hi_o[3])
         );
  OAI211V2_8TH40 U164 ( .A1(n32), .A2(n37), .B(n153), .C(n154), .ZN(hi_o[2])
         );
  OAI211V2_8TH40 U165 ( .A1(n190), .A2(n37), .B(n191), .C(n192), .ZN(hi_o[20])
         );
  OAI211V2_8TH40 U166 ( .A1(n33), .A2(n37), .B(n194), .C(n195), .ZN(hi_o[1])
         );
  OAI211V2_8TH40 U167 ( .A1(n197), .A2(n37), .B(n198), .C(n199), .ZN(hi_o[19])
         );
  OAI211V2_8TH40 U168 ( .A1(n22), .A2(n37), .B(n201), .C(n202), .ZN(hi_o[18])
         );
  OAI211V2_8TH40 U169 ( .A1(n23), .A2(n37), .B(n204), .C(n205), .ZN(hi_o[17])
         );
  OAI211V2_8TH40 U170 ( .A1(n24), .A2(n37), .B(n207), .C(n208), .ZN(hi_o[16])
         );
  OAI211V2_8TH40 U171 ( .A1(n210), .A2(n37), .B(n211), .C(n212), .ZN(hi_o[15])
         );
  OAI211V2_8TH40 U172 ( .A1(n214), .A2(n37), .B(n215), .C(n216), .ZN(hi_o[14])
         );
  OAI211V2_8TH40 U173 ( .A1(n25), .A2(n37), .B(n218), .C(n219), .ZN(hi_o[13])
         );
  OAI211V2_8TH40 U174 ( .A1(n221), .A2(n37), .B(n222), .C(n223), .ZN(hi_o[12])
         );
  OAI211V2_8TH40 U175 ( .A1(n26), .A2(n37), .B(n225), .C(n226), .ZN(hi_o[11])
         );
  OAI211V2_8TH40 U176 ( .A1(n27), .A2(n37), .B(n228), .C(n229), .ZN(hi_o[10])
         );
  OAI211V2_8TH40 U177 ( .A1(n231), .A2(n37), .B(n232), .C(n233), .ZN(hi_o[0])
         );
  OR2V4_8TH40 U178 ( .A1(maddmsub_stall_req), .A2(div_start), .Z(stall_req) );
  AOI22V2_8TH40 U179 ( .A1(div_res[9]), .A2(n40), .B1(mul_res_tmp1[9]), .B2(n3), .ZN(n39) );
  AOI22V2_8TH40 U180 ( .A1(div_res[8]), .A2(n40), .B1(mul_res_tmp1[8]), .B2(n3), .ZN(n44) );
  AOI22V2_8TH40 U181 ( .A1(div_res[7]), .A2(n40), .B1(mul_res_tmp1[7]), .B2(n3), .ZN(n46) );
  AOI22V2_8TH40 U182 ( .A1(div_res[6]), .A2(n40), .B1(mul_res_tmp1[6]), .B2(n3), .ZN(n48) );
  AOI22V2_8TH40 U183 ( .A1(div_res[5]), .A2(n40), .B1(mul_res_tmp1[5]), .B2(n3), .ZN(n50) );
  AOI22V2_8TH40 U184 ( .A1(div_res[4]), .A2(n40), .B1(mul_res_tmp1[4]), .B2(n3), .ZN(n52) );
  AOI22V2_8TH40 U185 ( .A1(div_res[3]), .A2(n40), .B1(mul_res_tmp1[3]), .B2(n3), .ZN(n54) );
  AOI22V2_8TH40 U186 ( .A1(div_res[31]), .A2(n40), .B1(mul_res_tmp1[31]), .B2(
        n3), .ZN(n56) );
  AOI22V2_8TH40 U187 ( .A1(div_res[30]), .A2(n40), .B1(mul_res_tmp1[30]), .B2(
        n3), .ZN(n58) );
  AOI22V2_8TH40 U188 ( .A1(div_res[2]), .A2(n40), .B1(mul_res_tmp1[2]), .B2(n3), .ZN(n60) );
  AOI22V2_8TH40 U189 ( .A1(div_res[29]), .A2(n40), .B1(mul_res_tmp1[29]), .B2(
        n3), .ZN(n62) );
  AOI22V2_8TH40 U190 ( .A1(div_res[28]), .A2(n40), .B1(mul_res_tmp1[28]), .B2(
        n3), .ZN(n64) );
  AOI22V2_8TH40 U191 ( .A1(div_res[27]), .A2(n40), .B1(mul_res_tmp1[27]), .B2(
        n3), .ZN(n66) );
  AOI22V2_8TH40 U192 ( .A1(div_res[26]), .A2(n40), .B1(mul_res_tmp1[26]), .B2(
        n3), .ZN(n68) );
  AOI22V2_8TH40 U193 ( .A1(div_res[25]), .A2(n40), .B1(mul_res_tmp1[25]), .B2(
        n3), .ZN(n70) );
  AOI22V2_8TH40 U194 ( .A1(div_res[24]), .A2(n40), .B1(mul_res_tmp1[24]), .B2(
        n3), .ZN(n72) );
  AOI22V2_8TH40 U195 ( .A1(div_res[23]), .A2(n40), .B1(mul_res_tmp1[23]), .B2(
        n3), .ZN(n74) );
  AOI22V2_8TH40 U196 ( .A1(div_res[22]), .A2(n40), .B1(mul_res_tmp1[22]), .B2(
        n3), .ZN(n76) );
  AOI22V2_8TH40 U197 ( .A1(div_res[21]), .A2(n40), .B1(mul_res_tmp1[21]), .B2(
        n3), .ZN(n78) );
  AOI22V2_8TH40 U198 ( .A1(div_res[20]), .A2(n40), .B1(mul_res_tmp1[20]), .B2(
        n3), .ZN(n80) );
  AOI22V2_8TH40 U199 ( .A1(div_res[1]), .A2(n40), .B1(mul_res_tmp1[1]), .B2(n3), .ZN(n82) );
  AOI22V2_8TH40 U200 ( .A1(div_res[19]), .A2(n40), .B1(mul_res_tmp1[19]), .B2(
        n3), .ZN(n84) );
  AOI22V2_8TH40 U201 ( .A1(div_res[18]), .A2(n40), .B1(mul_res_tmp1[18]), .B2(
        n3), .ZN(n86) );
  AOI22V2_8TH40 U202 ( .A1(div_res[17]), .A2(n40), .B1(mul_res_tmp1[17]), .B2(
        n3), .ZN(n88) );
  AOI22V2_8TH40 U203 ( .A1(div_res[16]), .A2(n40), .B1(mul_res_tmp1[16]), .B2(
        n3), .ZN(n90) );
  AOI22V2_8TH40 U204 ( .A1(div_res[15]), .A2(n40), .B1(mul_res_tmp1[15]), .B2(
        n3), .ZN(n92) );
  AOI22V2_8TH40 U205 ( .A1(div_res[14]), .A2(n40), .B1(mul_res_tmp1[14]), .B2(
        n3), .ZN(n94) );
  AOI22V2_8TH40 U206 ( .A1(div_res[13]), .A2(n40), .B1(mul_res_tmp1[13]), .B2(
        n3), .ZN(n96) );
  AOI22V2_8TH40 U207 ( .A1(div_res[12]), .A2(n40), .B1(mul_res_tmp1[12]), .B2(
        n3), .ZN(n98) );
  AOI22V2_8TH40 U208 ( .A1(div_res[11]), .A2(n40), .B1(mul_res_tmp1[11]), .B2(
        n3), .ZN(n100) );
  AOI22V2_8TH40 U209 ( .A1(div_res[10]), .A2(n40), .B1(mul_res_tmp1[10]), .B2(
        n3), .ZN(n102) );
  AOI22V2_8TH40 U210 ( .A1(div_res[0]), .A2(n40), .B1(mul_res_tmp1[0]), .B2(n3), .ZN(n104) );
  AOI22V2_8TH40 U211 ( .A1(div_res[41]), .A2(n40), .B1(mul_res_tmp1[41]), .B2(
        n3), .ZN(n123) );
  AOI22V2_8TH40 U212 ( .A1(div_res[40]), .A2(n40), .B1(mul_res_tmp1[40]), .B2(
        n3), .ZN(n126) );
  AOI22V2_8TH40 U213 ( .A1(div_res[39]), .A2(n40), .B1(mul_res_tmp1[39]), .B2(
        n3), .ZN(n130) );
  AOI22V2_8TH40 U214 ( .A1(div_res[38]), .A2(n40), .B1(mul_res_tmp1[38]), .B2(
        n3), .ZN(n133) );
  AOI22V2_8TH40 U215 ( .A1(div_res[37]), .A2(n40), .B1(mul_res_tmp1[37]), .B2(
        n3), .ZN(n137) );
  AOI22V2_8TH40 U216 ( .A1(div_res[36]), .A2(n40), .B1(mul_res_tmp1[36]), .B2(
        n3), .ZN(n140) );
  AOI22V2_8TH40 U217 ( .A1(div_res[35]), .A2(n40), .B1(mul_res_tmp1[35]), .B2(
        n3), .ZN(n144) );
  AOI22V2_8TH40 U218 ( .A1(div_res[34]), .A2(n40), .B1(mul_res_tmp1[34]), .B2(
        n3), .ZN(n154) );
  AOI22V2_8TH40 U219 ( .A1(div_res[52]), .A2(n40), .B1(mul_res_tmp1[52]), .B2(
        n3), .ZN(n192) );
  AOI22V2_8TH40 U220 ( .A1(div_res[33]), .A2(n40), .B1(mul_res_tmp1[33]), .B2(
        n3), .ZN(n195) );
  AOI22V2_8TH40 U221 ( .A1(div_res[51]), .A2(n40), .B1(mul_res_tmp1[51]), .B2(
        n3), .ZN(n199) );
  AOI22V2_8TH40 U222 ( .A1(div_res[50]), .A2(n40), .B1(mul_res_tmp1[50]), .B2(
        n3), .ZN(n202) );
  AOI22V2_8TH40 U223 ( .A1(div_res[49]), .A2(n40), .B1(mul_res_tmp1[49]), .B2(
        n3), .ZN(n205) );
  AOI22V2_8TH40 U224 ( .A1(div_res[48]), .A2(n40), .B1(mul_res_tmp1[48]), .B2(
        n3), .ZN(n208) );
  AOI22V2_8TH40 U225 ( .A1(div_res[47]), .A2(n40), .B1(mul_res_tmp1[47]), .B2(
        n3), .ZN(n212) );
  AOI22V2_8TH40 U226 ( .A1(div_res[46]), .A2(n40), .B1(mul_res_tmp1[46]), .B2(
        n3), .ZN(n216) );
  AOI22V2_8TH40 U227 ( .A1(div_res[45]), .A2(n40), .B1(mul_res_tmp1[45]), .B2(
        n3), .ZN(n219) );
  AOI22V2_8TH40 U228 ( .A1(div_res[44]), .A2(n40), .B1(mul_res_tmp1[44]), .B2(
        n3), .ZN(n223) );
  AOI22V2_8TH40 U229 ( .A1(div_res[43]), .A2(n40), .B1(mul_res_tmp1[43]), .B2(
        n3), .ZN(n226) );
  AOI22V2_8TH40 U230 ( .A1(div_res[42]), .A2(n40), .B1(mul_res_tmp1[42]), .B2(
        n3), .ZN(n229) );
  AOI22V2_8TH40 U231 ( .A1(div_res[32]), .A2(n40), .B1(mul_res_tmp1[32]), .B2(
        n3), .ZN(n233) );
  AOAOI2111V4_8TH40 U232 ( .A1(n745), .A2(inst_type[1]), .B(n755), .C(n802), 
        .D(n835), .ZN(n827) );
  AOA211V4_8TH40 U233 ( .A1(n234), .A2(n826), .B(n836), .C(n830), .Z(n835) );
  INOR2V2_8TH40 U234 ( .A1(n35), .B1(n1015), .ZN(n36) );
  INOR2V2_8TH40 U235 ( .A1(n35), .B1(n1042), .ZN(n34) );
  AOI222V2_8TH40 U236 ( .A1(mem_cp0_wdata[30]), .A2(n250), .B1(n251), .B2(n951), .C1(N1869), .C2(n252), .ZN(n420) );
  AOI222V2_8TH40 U237 ( .A1(mem_cp0_wdata[28]), .A2(n250), .B1(n251), .B2(n953), .C1(N1867), .C2(n252), .ZN(n484) );
  AOI222V2_8TH40 U238 ( .A1(mem_cp0_wdata[6]), .A2(n250), .B1(n251), .B2(n975), 
        .C1(N1845), .C2(n252), .ZN(n295) );
  AOI222V2_8TH40 U239 ( .A1(mem_cp0_wdata[13]), .A2(n250), .B1(n251), .B2(n968), .C1(N1852), .C2(n252), .ZN(n693) );
  AOI22V2_8TH40 U240 ( .A1(mul_res_tmp[44]), .A2(n843), .B1(N647), .B2(n844), 
        .ZN(n224) );
  AOI22V2_8TH40 U241 ( .A1(mul_res_tmp[45]), .A2(n843), .B1(N648), .B2(n844), 
        .ZN(n220) );
  AOI22V2_8TH40 U242 ( .A1(mul_res_tmp[4]), .A2(n843), .B1(N607), .B2(n844), 
        .ZN(n362) );
  AOI22V2_8TH40 U243 ( .A1(mul_res_tmp[5]), .A2(n843), .B1(N608), .B2(n844), 
        .ZN(n330) );
  AOI22V2_8TH40 U244 ( .A1(mul_res_tmp[6]), .A2(n843), .B1(N609), .B2(n844), 
        .ZN(n301) );
  AOI22V2_8TH40 U245 ( .A1(mul_res_tmp[7]), .A2(n843), .B1(N610), .B2(n844), 
        .ZN(n287) );
  AOI22V2_8TH40 U246 ( .A1(mul_res_tmp[8]), .A2(n843), .B1(N611), .B2(n844), 
        .ZN(n277) );
  AOI22V2_8TH40 U247 ( .A1(mul_res_tmp[9]), .A2(n843), .B1(N612), .B2(n844), 
        .ZN(n253) );
  AOI22V2_8TH40 U248 ( .A1(mul_res_tmp[10]), .A2(n843), .B1(N613), .B2(n844), 
        .ZN(n728) );
  AOI22V2_8TH40 U249 ( .A1(mul_res_tmp[12]), .A2(n843), .B1(N615), .B2(n844), 
        .ZN(n711) );
  AOI22V2_8TH40 U250 ( .A1(mul_res_tmp[13]), .A2(n843), .B1(N616), .B2(n844), 
        .ZN(n697) );
  AOI22V2_8TH40 U251 ( .A1(mul_res_tmp[14]), .A2(n843), .B1(N617), .B2(n844), 
        .ZN(n690) );
  AOI22V2_8TH40 U252 ( .A1(mul_res_tmp[15]), .A2(n843), .B1(N618), .B2(n844), 
        .ZN(n675) );
  AOI22V2_8TH40 U253 ( .A1(mul_res_tmp[20]), .A2(n843), .B1(N623), .B2(n844), 
        .ZN(n584) );
  AOI22V2_8TH40 U254 ( .A1(mul_res_tmp[21]), .A2(n843), .B1(N624), .B2(n844), 
        .ZN(n568) );
  AOI22V2_8TH40 U255 ( .A1(mul_res_tmp[22]), .A2(n843), .B1(N625), .B2(n844), 
        .ZN(n562) );
  AOI22V2_8TH40 U256 ( .A1(mul_res_tmp[24]), .A2(n843), .B1(N627), .B2(n844), 
        .ZN(n540) );
  AOI22V2_8TH40 U257 ( .A1(mul_res_tmp[25]), .A2(n843), .B1(N628), .B2(n844), 
        .ZN(n527) );
  AOI22V2_8TH40 U258 ( .A1(mul_res_tmp[26]), .A2(n843), .B1(N629), .B2(n844), 
        .ZN(n515) );
  AOI22V2_8TH40 U259 ( .A1(mul_res_tmp[27]), .A2(n843), .B1(N630), .B2(n844), 
        .ZN(n504) );
  AOI22V2_8TH40 U260 ( .A1(mul_res_tmp[28]), .A2(n843), .B1(N631), .B2(n844), 
        .ZN(n488) );
  AOI22V2_8TH40 U261 ( .A1(mul_res_tmp[29]), .A2(n843), .B1(N632), .B2(n844), 
        .ZN(n481) );
  AOI22V2_8TH40 U262 ( .A1(mul_res_tmp[46]), .A2(n843), .B1(N649), .B2(n844), 
        .ZN(n217) );
  AOI22V2_8TH40 U263 ( .A1(mul_res_tmp[47]), .A2(n843), .B1(N650), .B2(n844), 
        .ZN(n213) );
  AOI22V2_8TH40 U264 ( .A1(mul_res_tmp[48]), .A2(n843), .B1(N651), .B2(n844), 
        .ZN(n209) );
  AOI22V2_8TH40 U265 ( .A1(mul_res_tmp[49]), .A2(n843), .B1(N652), .B2(n844), 
        .ZN(n206) );
  AOI22V2_8TH40 U266 ( .A1(mul_res_tmp[50]), .A2(n843), .B1(N653), .B2(n844), 
        .ZN(n203) );
  AOI22V2_8TH40 U267 ( .A1(mul_res_tmp[51]), .A2(n843), .B1(N654), .B2(n844), 
        .ZN(n200) );
  AOI22V2_8TH40 U268 ( .A1(mul_res_tmp[52]), .A2(n843), .B1(N655), .B2(n844), 
        .ZN(n193) );
  AOI22V2_8TH40 U269 ( .A1(mul_res_tmp[53]), .A2(n843), .B1(N656), .B2(n844), 
        .ZN(n189) );
  AOI22V2_8TH40 U270 ( .A1(mul_res_tmp[54]), .A2(n843), .B1(N657), .B2(n844), 
        .ZN(n186) );
  AOI22V2_8TH40 U271 ( .A1(mul_res_tmp[55]), .A2(n843), .B1(N658), .B2(n844), 
        .ZN(n182) );
  AOI22V2_8TH40 U272 ( .A1(mul_res_tmp[56]), .A2(n843), .B1(N659), .B2(n844), 
        .ZN(n178) );
  AOI22V2_8TH40 U273 ( .A1(mul_res_tmp[57]), .A2(n843), .B1(N660), .B2(n844), 
        .ZN(n174) );
  AOI22V2_8TH40 U274 ( .A1(mul_res_tmp[58]), .A2(n843), .B1(N661), .B2(n844), 
        .ZN(n170) );
  AOI22V2_8TH40 U275 ( .A1(mul_res_tmp[59]), .A2(n843), .B1(N662), .B2(n844), 
        .ZN(n166) );
  AOI22V2_8TH40 U276 ( .A1(mul_res_tmp[60]), .A2(n843), .B1(N663), .B2(n844), 
        .ZN(n162) );
  AOI22V2_8TH40 U277 ( .A1(mul_res_tmp[61]), .A2(n843), .B1(N664), .B2(n844), 
        .ZN(n159) );
  AOI22V2_8TH40 U278 ( .A1(mul_res_tmp[62]), .A2(n843), .B1(N665), .B2(n844), 
        .ZN(n152) );
  NOR3V2_8TH40 U279 ( .A1(N1875), .A2(n664), .A3(n17), .ZN(n688) );
  AOI22V2_8TH40 U280 ( .A1(n251), .A2(n1013), .B1(N1839), .B2(n252), .ZN(n733)
         );
  AOI22V2_8TH40 U281 ( .A1(n251), .A2(n950), .B1(N1870), .B2(n252), .ZN(n406)
         );
  AOI22V2_8TH40 U282 ( .A1(n251), .A2(n978), .B1(N1842), .B2(n252), .ZN(n368)
         );
  NAND2V2_8TH40 U283 ( .A1(n269), .A2(n756), .ZN(n263) );
  INV2_8TH40 U284 ( .I(N951), .ZN(n906) );
  INV2_8TH40 U285 ( .I(N952), .ZN(n905) );
  INV2_8TH40 U286 ( .I(N953), .ZN(n904) );
  INV2_8TH40 U287 ( .I(N954), .ZN(n903) );
  INV2_8TH40 U288 ( .I(N955), .ZN(n902) );
  INV2_8TH40 U289 ( .I(N956), .ZN(n901) );
  INV2_8TH40 U290 ( .I(N957), .ZN(n900) );
  INV2_8TH40 U291 ( .I(N958), .ZN(n899) );
  INV2_8TH40 U292 ( .I(N959), .ZN(n898) );
  INV2_8TH40 U293 ( .I(N960), .ZN(n897) );
  INV2_8TH40 U294 ( .I(N961), .ZN(n896) );
  INV2_8TH40 U295 ( .I(N962), .ZN(n895) );
  INV2_8TH40 U296 ( .I(N963), .ZN(n894) );
  INV2_8TH40 U297 ( .I(N964), .ZN(n893) );
  INV2_8TH40 U298 ( .I(N965), .ZN(n892) );
  INV2_8TH40 U299 ( .I(N966), .ZN(n891) );
  INV2_8TH40 U300 ( .I(N967), .ZN(n890) );
  INV2_8TH40 U301 ( .I(N968), .ZN(n889) );
  INV2_8TH40 U302 ( .I(N969), .ZN(n888) );
  INV2_8TH40 U303 ( .I(N970), .ZN(n887) );
  INV2_8TH40 U304 ( .I(N971), .ZN(n886) );
  OAI22V2_8TH40 U305 ( .A1(n562), .A2(n838), .B1(n885), .B2(n842), .ZN(N1370)
         );
  INV2_8TH40 U306 ( .I(N972), .ZN(n885) );
  OAI22V2_8TH40 U307 ( .A1(n546), .A2(n838), .B1(n884), .B2(n842), .ZN(N1371)
         );
  INV2_8TH40 U308 ( .I(N973), .ZN(n884) );
  OAI22V2_8TH40 U309 ( .A1(n540), .A2(n838), .B1(n883), .B2(n842), .ZN(N1372)
         );
  INV2_8TH40 U310 ( .I(N974), .ZN(n883) );
  OAI22V2_8TH40 U311 ( .A1(n527), .A2(n838), .B1(n882), .B2(n842), .ZN(N1373)
         );
  INV2_8TH40 U312 ( .I(N975), .ZN(n882) );
  OAI22V2_8TH40 U313 ( .A1(n515), .A2(n838), .B1(n881), .B2(n842), .ZN(N1374)
         );
  INV2_8TH40 U314 ( .I(N976), .ZN(n881) );
  OAI22V2_8TH40 U315 ( .A1(n504), .A2(n838), .B1(n880), .B2(n842), .ZN(N1375)
         );
  INV2_8TH40 U316 ( .I(N977), .ZN(n880) );
  OAI22V2_8TH40 U317 ( .A1(n488), .A2(n838), .B1(n879), .B2(n842), .ZN(N1376)
         );
  INV2_8TH40 U318 ( .I(N978), .ZN(n879) );
  OAI22V2_8TH40 U319 ( .A1(n481), .A2(n838), .B1(n878), .B2(n842), .ZN(N1377)
         );
  INV2_8TH40 U320 ( .I(N979), .ZN(n878) );
  OAI22V2_8TH40 U321 ( .A1(n425), .A2(n838), .B1(n877), .B2(n842), .ZN(N1378)
         );
  INV2_8TH40 U322 ( .I(N980), .ZN(n877) );
  OAI22V2_8TH40 U323 ( .A1(n417), .A2(n838), .B1(n876), .B2(n842), .ZN(N1379)
         );
  INV2_8TH40 U324 ( .I(N981), .ZN(n876) );
  OAI22V2_8TH40 U325 ( .A1(n237), .A2(n838), .B1(n875), .B2(n842), .ZN(N1380)
         );
  INV2_8TH40 U326 ( .I(N982), .ZN(n875) );
  OAI22V2_8TH40 U327 ( .A1(n196), .A2(n838), .B1(n874), .B2(n842), .ZN(N1381)
         );
  INV2_8TH40 U328 ( .I(N983), .ZN(n874) );
  OAI22V2_8TH40 U329 ( .A1(n155), .A2(n838), .B1(n873), .B2(n842), .ZN(N1382)
         );
  INV2_8TH40 U330 ( .I(N984), .ZN(n873) );
  OAI22V2_8TH40 U331 ( .A1(n145), .A2(n838), .B1(n872), .B2(n842), .ZN(N1383)
         );
  INV2_8TH40 U332 ( .I(N985), .ZN(n872) );
  OAI22V2_8TH40 U333 ( .A1(n141), .A2(n838), .B1(n871), .B2(n842), .ZN(N1384)
         );
  INV2_8TH40 U334 ( .I(N986), .ZN(n871) );
  OAI22V2_8TH40 U335 ( .A1(n138), .A2(n838), .B1(n870), .B2(n842), .ZN(N1385)
         );
  INV2_8TH40 U336 ( .I(N987), .ZN(n870) );
  OAI22V2_8TH40 U337 ( .A1(n134), .A2(n838), .B1(n869), .B2(n842), .ZN(N1386)
         );
  INV2_8TH40 U338 ( .I(N988), .ZN(n869) );
  OAI22V2_8TH40 U339 ( .A1(n131), .A2(n838), .B1(n868), .B2(n842), .ZN(N1387)
         );
  INV2_8TH40 U340 ( .I(N989), .ZN(n868) );
  OAI22V2_8TH40 U341 ( .A1(n127), .A2(n838), .B1(n867), .B2(n842), .ZN(N1388)
         );
  INV2_8TH40 U342 ( .I(N990), .ZN(n867) );
  OAI22V2_8TH40 U343 ( .A1(n124), .A2(n838), .B1(n866), .B2(n842), .ZN(N1389)
         );
  INV2_8TH40 U344 ( .I(N991), .ZN(n866) );
  OAI22V2_8TH40 U345 ( .A1(n230), .A2(n838), .B1(n865), .B2(n842), .ZN(N1390)
         );
  INV2_8TH40 U346 ( .I(N992), .ZN(n865) );
  OAI22V2_8TH40 U347 ( .A1(n227), .A2(n838), .B1(n864), .B2(n842), .ZN(N1391)
         );
  INV2_8TH40 U348 ( .I(N993), .ZN(n864) );
  OAI22V2_8TH40 U349 ( .A1(n224), .A2(n838), .B1(n863), .B2(n842), .ZN(N1392)
         );
  INV2_8TH40 U350 ( .I(N994), .ZN(n863) );
  OAI22V2_8TH40 U351 ( .A1(n220), .A2(n838), .B1(n862), .B2(n842), .ZN(N1393)
         );
  INV2_8TH40 U352 ( .I(N995), .ZN(n862) );
  OAI22V2_8TH40 U353 ( .A1(n217), .A2(n838), .B1(n861), .B2(n842), .ZN(N1394)
         );
  INV2_8TH40 U354 ( .I(N996), .ZN(n861) );
  OAI22V2_8TH40 U355 ( .A1(n213), .A2(n838), .B1(n860), .B2(n842), .ZN(N1395)
         );
  INV2_8TH40 U356 ( .I(N997), .ZN(n860) );
  OAI22V2_8TH40 U357 ( .A1(n209), .A2(n838), .B1(n859), .B2(n842), .ZN(N1396)
         );
  INV2_8TH40 U358 ( .I(N998), .ZN(n859) );
  OAI22V2_8TH40 U359 ( .A1(n206), .A2(n838), .B1(n858), .B2(n842), .ZN(N1397)
         );
  INV2_8TH40 U360 ( .I(N999), .ZN(n858) );
  OAI22V2_8TH40 U361 ( .A1(n203), .A2(n838), .B1(n857), .B2(n842), .ZN(N1398)
         );
  INV2_8TH40 U362 ( .I(N1000), .ZN(n857) );
  OAI22V2_8TH40 U363 ( .A1(n200), .A2(n838), .B1(n856), .B2(n842), .ZN(N1399)
         );
  INV2_8TH40 U364 ( .I(N1001), .ZN(n856) );
  OAI22V2_8TH40 U365 ( .A1(n193), .A2(n838), .B1(n855), .B2(n842), .ZN(N1400)
         );
  INV2_8TH40 U366 ( .I(N1002), .ZN(n855) );
  OAI22V2_8TH40 U367 ( .A1(n189), .A2(n838), .B1(n854), .B2(n842), .ZN(N1401)
         );
  INV2_8TH40 U368 ( .I(N1003), .ZN(n854) );
  OAI22V2_8TH40 U369 ( .A1(n186), .A2(n838), .B1(n853), .B2(n842), .ZN(N1402)
         );
  INV2_8TH40 U370 ( .I(N1004), .ZN(n853) );
  OAI22V2_8TH40 U371 ( .A1(n182), .A2(n838), .B1(n852), .B2(n842), .ZN(N1403)
         );
  INV2_8TH40 U372 ( .I(N1005), .ZN(n852) );
  OAI22V2_8TH40 U373 ( .A1(n178), .A2(n838), .B1(n851), .B2(n842), .ZN(N1404)
         );
  INV2_8TH40 U374 ( .I(N1006), .ZN(n851) );
  OAI22V2_8TH40 U375 ( .A1(n174), .A2(n838), .B1(n850), .B2(n842), .ZN(N1405)
         );
  INV2_8TH40 U376 ( .I(N1007), .ZN(n850) );
  OAI22V2_8TH40 U377 ( .A1(n170), .A2(n838), .B1(n849), .B2(n842), .ZN(N1406)
         );
  INV2_8TH40 U378 ( .I(N1008), .ZN(n849) );
  OAI22V2_8TH40 U379 ( .A1(n166), .A2(n838), .B1(n848), .B2(n842), .ZN(N1407)
         );
  INV2_8TH40 U380 ( .I(N1009), .ZN(n848) );
  OAI22V2_8TH40 U381 ( .A1(n162), .A2(n838), .B1(n847), .B2(n842), .ZN(N1408)
         );
  INV2_8TH40 U382 ( .I(N1010), .ZN(n847) );
  OAI22V2_8TH40 U383 ( .A1(n159), .A2(n838), .B1(n846), .B2(n842), .ZN(N1409)
         );
  INV2_8TH40 U384 ( .I(N1011), .ZN(n846) );
  OAI22V2_8TH40 U385 ( .A1(n152), .A2(n838), .B1(n845), .B2(n842), .ZN(N1410)
         );
  INV2_8TH40 U386 ( .I(N1012), .ZN(n845) );
  INV2_8TH40 U387 ( .I(N1013), .ZN(n841) );
  OAI22V2_8TH40 U388 ( .A1(n907), .A2(n239), .B1(n840), .B2(n807), .ZN(n35) );
  AOI31V2_8TH40 U389 ( .A1(n238), .A2(n764), .A3(n742), .B(n908), .ZN(n907) );
  AOI22V2_8TH40 U390 ( .A1(N1840), .A2(n252), .B1(mem_cp0_wdata[1]), .B2(n250), 
        .ZN(n592) );
  AOI22V2_8TH40 U391 ( .A1(N1841), .A2(n252), .B1(mem_cp0_wdata[2]), .B2(n250), 
        .ZN(n437) );
  OAI32V2_8TH40 U392 ( .A1(n791), .A2(n762), .A3(n792), .B1(n276), .B2(n299), 
        .ZN(n780) );
  NAND4V2_8TH40 U393 ( .A1(n573), .A2(n574), .A3(n575), .A4(n576), .ZN(
        exe_result_o[20]) );
  I2NOR3V2_8TH40 U394 ( .A1(n577), .A2(n578), .B(n579), .ZN(n576) );
  MAOI22V2_8TH40 U395 ( .A1(sum_res[20]), .A2(n244), .B1(n548), .B2(n353), 
        .ZN(n574) );
  AOI222V2_8TH40 U396 ( .A1(n288), .A2(lo[20]), .B1(N1859), .B2(n252), .C1(
        mem_cp0_wdata[20]), .C2(n250), .ZN(n575) );
  NAND4V2_8TH40 U397 ( .A1(n551), .A2(n552), .A3(n553), .A4(n554), .ZN(
        exe_result_o[22]) );
  I2NOR3V2_8TH40 U398 ( .A1(n555), .A2(n556), .B(n557), .ZN(n554) );
  MAOI22V2_8TH40 U399 ( .A1(sum_res[22]), .A2(n244), .B1(n548), .B2(n298), 
        .ZN(n552) );
  AOI222V2_8TH40 U400 ( .A1(n288), .A2(lo[22]), .B1(N1861), .B2(n252), .C1(
        mem_cp0_wdata[22]), .C2(n250), .ZN(n553) );
  NAND4V2_8TH40 U401 ( .A1(n528), .A2(n529), .A3(n530), .A4(n531), .ZN(
        exe_result_o[24]) );
  I2NOR3V2_8TH40 U402 ( .A1(n532), .A2(n533), .B(n534), .ZN(n531) );
  AOI22V2_8TH40 U403 ( .A1(n416), .A2(n539), .B1(sum_res[24]), .B2(n244), .ZN(
        n529) );
  AOI222V2_8TH40 U404 ( .A1(n288), .A2(lo[24]), .B1(N1863), .B2(n252), .C1(
        mem_cp0_wdata[24]), .C2(n250), .ZN(n530) );
  NAND4V2_8TH40 U405 ( .A1(n516), .A2(n517), .A3(n518), .A4(n519), .ZN(
        exe_result_o[25]) );
  I2NOR3V2_8TH40 U406 ( .A1(n520), .A2(n521), .B(n522), .ZN(n519) );
  AOI22V2_8TH40 U407 ( .A1(n416), .A2(n526), .B1(sum_res[25]), .B2(n244), .ZN(
        n517) );
  AOI222V2_8TH40 U408 ( .A1(n288), .A2(lo[25]), .B1(N1864), .B2(n252), .C1(
        mem_cp0_wdata[25]), .C2(n250), .ZN(n518) );
  NAND4V2_8TH40 U409 ( .A1(n505), .A2(n506), .A3(n507), .A4(n508), .ZN(
        exe_result_o[26]) );
  I2NOR3V2_8TH40 U410 ( .A1(n509), .A2(n510), .B(n511), .ZN(n508) );
  AOI22V2_8TH40 U411 ( .A1(n441), .A2(n416), .B1(sum_res[26]), .B2(n244), .ZN(
        n506) );
  AOI222V2_8TH40 U412 ( .A1(n288), .A2(lo[26]), .B1(N1865), .B2(n252), .C1(
        mem_cp0_wdata[26]), .C2(n250), .ZN(n507) );
  NAND4V2_8TH40 U413 ( .A1(n493), .A2(n494), .A3(n495), .A4(n496), .ZN(
        exe_result_o[27]) );
  I2NOR3V2_8TH40 U414 ( .A1(n497), .A2(n498), .B(n499), .ZN(n496) );
  AOI22V2_8TH40 U415 ( .A1(n416), .A2(n503), .B1(sum_res[27]), .B2(n244), .ZN(
        n494) );
  AOI222V2_8TH40 U416 ( .A1(n288), .A2(lo[27]), .B1(N1866), .B2(n252), .C1(
        mem_cp0_wdata[27]), .C2(n250), .ZN(n495) );
  NAND4V2_8TH40 U417 ( .A1(n469), .A2(n470), .A3(n471), .A4(n472), .ZN(
        exe_result_o[29]) );
  I2NOR3V2_8TH40 U418 ( .A1(n473), .A2(n474), .B(n475), .ZN(n472) );
  AOI22V2_8TH40 U419 ( .A1(n416), .A2(n329), .B1(sum_res[29]), .B2(n244), .ZN(
        n470) );
  AOI222V2_8TH40 U420 ( .A1(n288), .A2(lo[29]), .B1(N1868), .B2(n252), .C1(
        mem_cp0_wdata[29]), .C2(n250), .ZN(n471) );
  NAND4V2_8TH40 U421 ( .A1(n306), .A2(n307), .A3(n308), .A4(n309), .ZN(
        exe_result_o[5]) );
  AOI22V2_8TH40 U422 ( .A1(n328), .A2(n329), .B1(sum_res[5]), .B2(n244), .ZN(
        n307) );
  I2NOR4V2_8TH40 U423 ( .A1(n310), .A2(n311), .B1(n312), .B2(n313), .ZN(n309)
         );
  AOI222V2_8TH40 U424 ( .A1(n288), .A2(lo[5]), .B1(N1844), .B2(n252), .C1(
        mem_cp0_wdata[5]), .C2(n250), .ZN(n308) );
  NAND4V2_8TH40 U425 ( .A1(n702), .A2(n703), .A3(n704), .A4(n705), .ZN(
        exe_result_o[12]) );
  I2NOR3V2_8TH40 U426 ( .A1(n706), .A2(n707), .B(n708), .ZN(n705) );
  AOI22V2_8TH40 U427 ( .A1(n688), .A2(n487), .B1(sum_res[12]), .B2(n244), .ZN(
        n703) );
  AOI222V2_8TH40 U428 ( .A1(n288), .A2(lo[12]), .B1(N1851), .B2(n252), .C1(
        mem_cp0_wdata[12]), .C2(n250), .ZN(n704) );
  NAND4V2_8TH40 U429 ( .A1(n679), .A2(n680), .A3(n681), .A4(n682), .ZN(
        exe_result_o[14]) );
  I2NOR3V2_8TH40 U430 ( .A1(n683), .A2(n684), .B(n685), .ZN(n682) );
  AOI22V2_8TH40 U431 ( .A1(n688), .A2(n423), .B1(sum_res[14]), .B2(n244), .ZN(
        n680) );
  AOI222V2_8TH40 U432 ( .A1(n288), .A2(lo[14]), .B1(N1853), .B2(n252), .C1(
        mem_cp0_wdata[14]), .C2(n250), .ZN(n681) );
  NAND4V2_8TH40 U433 ( .A1(n331), .A2(n332), .A3(n333), .A4(n334), .ZN(
        exe_result_o[4]) );
  AOI211V2_8TH40 U434 ( .A1(sum_res[4]), .A2(n244), .B(n342), .C(n343), .ZN(
        n333) );
  AOI22V2_8TH40 U435 ( .A1(N1843), .A2(n252), .B1(mem_cp0_wdata[4]), .B2(n250), 
        .ZN(n331) );
  INOR4V2_8TH40 U436 ( .A1(n335), .B1(n336), .B2(n337), .B3(n338), .ZN(n334)
         );
  AOI22V2_8TH40 U437 ( .A1(n820), .A2(n821), .B1(n817), .B2(n760), .ZN(n813)
         );
  I2NOR4V2_8TH40 U438 ( .A1(n235), .A2(n238), .B1(n239), .B2(inst_type[1]), 
        .ZN(n41) );
  NOR3V2_8TH40 U439 ( .A1(df_wbex_hilo_we), .A2(rst), .A3(df_memex_hilo_we), 
        .ZN(n261) );
  AOI21V2_8TH40 U440 ( .A1(n35), .A2(n414), .B(rst), .ZN(n843) );
  INAND3V2_8TH40 U441 ( .A1(n840), .B1(n759), .B2(n909), .ZN(n842) );
  NAND2V0_8TH40 U442 ( .A1(cycl_cnt_i[1]), .A2(n3), .ZN(N1413) );
  NAND4V2_8TH40 U443 ( .A1(n810), .A2(inst_type[6]), .A3(n742), .A4(n825), 
        .ZN(n824) );
  AND4V2_8TH40 U444 ( .A1(n742), .A2(inst_type[6]), .A3(n743), .A4(n744), .Z(
        n262) );
  INV2_8TH40 U445 ( .I(n801), .ZN(n244) );
  OAOAI2111V2_8TH40 U446 ( .A1(n802), .A2(n803), .B(n745), .C(n804), .D(n805), 
        .ZN(n801) );
  AOI222V2_8TH40 U447 ( .A1(mem_cp0_wdata[16]), .A2(n250), .B1(n251), .B2(n965), .C1(N1855), .C2(n252), .ZN(n661) );
  AOI222V2_8TH40 U448 ( .A1(mem_cp0_wdata[17]), .A2(n250), .B1(n251), .B2(n964), .C1(N1856), .C2(n252), .ZN(n651) );
  AOI222V2_8TH40 U449 ( .A1(mem_cp0_wdata[18]), .A2(n250), .B1(n251), .B2(n963), .C1(N1857), .C2(n252), .ZN(n640) );
  AOI222V2_8TH40 U450 ( .A1(mem_cp0_wdata[21]), .A2(n250), .B1(n251), .B2(n960), .C1(N1860), .C2(n252), .ZN(n565) );
  AOI221V2_8TH40 U451 ( .A1(link_addr[7]), .A2(n245), .B1(n251), .B2(n974), 
        .C(n286), .ZN(n285) );
  AOI221V2_8TH40 U452 ( .A1(link_addr[15]), .A2(n245), .B1(n251), .B2(n966), 
        .C(n674), .ZN(n673) );
  AOI221V2_8TH40 U453 ( .A1(n251), .A2(n962), .B1(N1858), .B2(n252), .C(n632), 
        .ZN(n631) );
  AO22V2_8TH40 U454 ( .A1(link_addr[19]), .A2(n245), .B1(sum_res[19]), .B2(
        n244), .Z(n632) );
  AOI221V2_8TH40 U455 ( .A1(n251), .A2(n958), .B1(N1862), .B2(n252), .C(n545), 
        .ZN(n544) );
  AO22V2_8TH40 U456 ( .A1(link_addr[23]), .A2(n245), .B1(sum_res[23]), .B2(
        n244), .Z(n545) );
  I2NOR4V2_8TH40 U457 ( .A1(n760), .A2(n761), .B1(n762), .B2(n763), .ZN(n754)
         );
  OAI221V2_8TH40 U458 ( .A1(n108), .A2(n258), .B1(n31), .B2(n257), .C(n341), 
        .ZN(n337) );
  AOI22V2_8TH40 U459 ( .A1(cp0_ex_rdata[4]), .A2(n254), .B1(wb_cp0_wdata[4]), 
        .B2(n255), .ZN(n341) );
  AOI222V2_8TH40 U460 ( .A1(wb_cp0_wdata[12]), .A2(n255), .B1(n289), .B2(n1000), .C1(cp0_ex_rdata[12]), .C2(n254), .ZN(n707) );
  AOI222V2_8TH40 U461 ( .A1(wb_cp0_wdata[14]), .A2(n255), .B1(n289), .B2(n998), 
        .C1(cp0_ex_rdata[14]), .C2(n254), .ZN(n684) );
  AOI222V2_8TH40 U462 ( .A1(wb_cp0_wdata[31]), .A2(n255), .B1(n266), .B2(n414), 
        .C1(cp0_ex_rdata[31]), .C2(n254), .ZN(n411) );
  I2NOR4V2_8TH40 U463 ( .A1(inst_class[1]), .A2(n811), .B1(inst_class[0]), 
        .B2(inst_class[2]), .ZN(n743) );
  OAI221V2_8TH40 U464 ( .A1(n393), .A2(n358), .B1(n394), .B2(n346), .C(n300), 
        .ZN(n336) );
  AOI211V2_8TH40 U465 ( .A1(n382), .A2(gpr1_data[7]), .B(n398), .C(n399), .ZN(
        n393) );
  AOI221V2_8TH40 U466 ( .A1(cp0_ex_rdata[1]), .A2(n254), .B1(wb_cp0_wdata[1]), 
        .B2(n255), .C(n589), .ZN(n587) );
  AOI221V2_8TH40 U467 ( .A1(cp0_ex_rdata[2]), .A2(n254), .B1(wb_cp0_wdata[2]), 
        .B2(n255), .C(n434), .ZN(n432) );
  AOI33V2_8TH40 U468 ( .A1(n790), .A2(n1040), .A3(gpr1_data[7]), .B1(n325), 
        .B2(n912), .B3(gpr1_data[1]), .ZN(n389) );
  MUX2V0_8TH40 U469 ( .I0(N60), .I1(gpr2_data[0]), .S(n827), .Z(
        com_gpr2_data[0]) );
  AOI211V2_8TH40 U470 ( .A1(n263), .A2(gpr1_data[3]), .B(n392), .C(n336), .ZN(
        n365) );
  MUX3V2_8TH40 U471 ( .I0(n265), .I1(n266), .I2(n404), .S0(gpr1_data[3]), .S1(
        gpr2_data[3]), .Z(n392) );
  NAND2V2_8TH40 U472 ( .A1(n405), .A2(n269), .ZN(n404) );
  OAI211V2_8TH40 U473 ( .A1(gpr1_data[16]), .A2(n350), .B(n619), .C(n620), 
        .ZN(n463) );
  OAOI211V2_8TH40 U474 ( .A1(n913), .A2(n912), .B(n325), .C(n621), .ZN(n620)
         );
  AOI22V2_8TH40 U475 ( .A1(wb_cp0_wdata[5]), .A2(n255), .B1(N1812), .B2(n262), 
        .ZN(n310) );
  OAI211V2_8TH40 U476 ( .A1(n1030), .A2(n359), .B(n603), .C(n604), .ZN(n449)
         );
  OAOI211V2_8TH40 U477 ( .A1(gpr1_data[0]), .A2(gpr1_data[1]), .B(n327), .C(
        n605), .ZN(n604) );
  OAOI211V2_8TH40 U478 ( .A1(gpr1_data[24]), .A2(gpr1_data[25]), .B(n607), .C(
        n608), .ZN(n603) );
  INAND4V2_8TH40 U479 ( .A1(n585), .B1(n586), .B2(n587), .B3(n588), .ZN(
        exe_result_o[1]) );
  MUX3V2_8TH40 U480 ( .I0(n316), .I1(n317), .I2(n590), .S0(gpr1_data[1]), .S1(
        gpr2_data[1]), .Z(n586) );
  NAND4V2_8TH40 U481 ( .A1(n592), .A2(n593), .A3(n594), .A4(n595), .ZN(n585)
         );
  AOI22V2_8TH40 U482 ( .A1(N1808), .A2(n262), .B1(n263), .B2(gpr1_data[1]), 
        .ZN(n588) );
  INAND4V2_8TH40 U483 ( .A1(n430), .B1(n431), .B2(n432), .B3(n433), .ZN(
        exe_result_o[2]) );
  MUX3V2_8TH40 U484 ( .I0(n316), .I1(n317), .I2(n435), .S0(gpr1_data[2]), .S1(
        gpr2_data[2]), .Z(n431) );
  NAND4V2_8TH40 U485 ( .A1(n437), .A2(n438), .A3(n439), .A4(n440), .ZN(n430)
         );
  AOI22V2_8TH40 U486 ( .A1(N1809), .A2(n262), .B1(n263), .B2(gpr1_data[2]), 
        .ZN(n433) );
  NAND4V2_8TH40 U487 ( .A1(n659), .A2(n660), .A3(n661), .A4(n662), .ZN(
        exe_result_o[16]) );
  AOI221V2_8TH40 U488 ( .A1(cp0_ex_rdata[16]), .A2(n254), .B1(wb_cp0_wdata[16]), .B2(n255), .C(n666), .ZN(n660) );
  AOI221V2_8TH40 U489 ( .A1(N1823), .A2(n262), .B1(n263), .B2(gpr1_data[16]), 
        .C(n667), .ZN(n659) );
  AOI221V2_8TH40 U490 ( .A1(sum_res[16]), .A2(n244), .B1(link_addr[16]), .B2(
        n245), .C(n663), .ZN(n662) );
  NAND4V2_8TH40 U491 ( .A1(n649), .A2(n650), .A3(n651), .A4(n652), .ZN(
        exe_result_o[17]) );
  AOI221V2_8TH40 U492 ( .A1(cp0_ex_rdata[17]), .A2(n254), .B1(wb_cp0_wdata[17]), .B2(n255), .C(n655), .ZN(n650) );
  AOI221V2_8TH40 U493 ( .A1(N1824), .A2(n262), .B1(n263), .B2(gpr1_data[17]), 
        .C(n656), .ZN(n649) );
  AOI221V2_8TH40 U494 ( .A1(sum_res[17]), .A2(n244), .B1(link_addr[17]), .B2(
        n245), .C(n653), .ZN(n652) );
  NAND4V2_8TH40 U495 ( .A1(n638), .A2(n639), .A3(n640), .A4(n641), .ZN(
        exe_result_o[18]) );
  AOI221V2_8TH40 U496 ( .A1(cp0_ex_rdata[18]), .A2(n254), .B1(wb_cp0_wdata[18]), .B2(n255), .C(n645), .ZN(n639) );
  AOI221V2_8TH40 U497 ( .A1(N1825), .A2(n262), .B1(n263), .B2(gpr1_data[18]), 
        .C(n646), .ZN(n638) );
  AOI221V2_8TH40 U498 ( .A1(sum_res[18]), .A2(n244), .B1(link_addr[18]), .B2(
        n245), .C(n642), .ZN(n641) );
  NAND4V2_8TH40 U499 ( .A1(n563), .A2(n564), .A3(n565), .A4(n566), .ZN(
        exe_result_o[21]) );
  AOI221V2_8TH40 U500 ( .A1(cp0_ex_rdata[21]), .A2(n254), .B1(wb_cp0_wdata[21]), .B2(n255), .C(n569), .ZN(n564) );
  AOI221V2_8TH40 U501 ( .A1(N1828), .A2(n262), .B1(n263), .B2(gpr1_data[21]), 
        .C(n570), .ZN(n563) );
  AOI221V2_8TH40 U502 ( .A1(sum_res[21]), .A2(n244), .B1(link_addr[21]), .B2(
        n245), .C(n567), .ZN(n566) );
  NAND4V2_8TH40 U503 ( .A1(n482), .A2(n483), .A3(n484), .A4(n485), .ZN(
        exe_result_o[28]) );
  AOI221V2_8TH40 U504 ( .A1(cp0_ex_rdata[28]), .A2(n254), .B1(wb_cp0_wdata[28]), .B2(n255), .C(n489), .ZN(n483) );
  AOI221V2_8TH40 U505 ( .A1(N1835), .A2(n262), .B1(n263), .B2(gpr1_data[28]), 
        .C(n490), .ZN(n482) );
  AOI221V2_8TH40 U506 ( .A1(sum_res[28]), .A2(n244), .B1(link_addr[28]), .B2(
        n245), .C(n486), .ZN(n485) );
  NAND4V2_8TH40 U507 ( .A1(n418), .A2(n419), .A3(n420), .A4(n421), .ZN(
        exe_result_o[30]) );
  AOI221V2_8TH40 U508 ( .A1(cp0_ex_rdata[30]), .A2(n254), .B1(wb_cp0_wdata[30]), .B2(n255), .C(n426), .ZN(n419) );
  AOI221V2_8TH40 U509 ( .A1(N1837), .A2(n262), .B1(n263), .B2(gpr1_data[30]), 
        .C(n427), .ZN(n418) );
  AOI221V2_8TH40 U510 ( .A1(sum_res[30]), .A2(n244), .B1(link_addr[30]), .B2(
        n245), .C(n422), .ZN(n421) );
  NAND4V2_8TH40 U511 ( .A1(n293), .A2(n294), .A3(n295), .A4(n296), .ZN(
        exe_result_o[6]) );
  AOI221V2_8TH40 U512 ( .A1(cp0_ex_rdata[6]), .A2(n254), .B1(wb_cp0_wdata[6]), 
        .B2(n255), .C(n302), .ZN(n294) );
  AOI221V2_8TH40 U513 ( .A1(N1813), .A2(n262), .B1(n263), .B2(gpr1_data[6]), 
        .C(n303), .ZN(n293) );
  AOI221V2_8TH40 U514 ( .A1(sum_res[6]), .A2(n244), .B1(link_addr[6]), .B2(
        n245), .C(n297), .ZN(n296) );
  NAND4V2_8TH40 U515 ( .A1(n271), .A2(n272), .A3(n273), .A4(n274), .ZN(
        exe_result_o[8]) );
  AOI221V2_8TH40 U516 ( .A1(cp0_ex_rdata[8]), .A2(n254), .B1(wb_cp0_wdata[8]), 
        .B2(n255), .C(n278), .ZN(n272) );
  AOI221V2_8TH40 U517 ( .A1(N1815), .A2(n262), .B1(n263), .B2(gpr1_data[8]), 
        .C(n279), .ZN(n271) );
  AOI221V2_8TH40 U518 ( .A1(sum_res[8]), .A2(n244), .B1(link_addr[8]), .B2(
        n245), .C(n275), .ZN(n274) );
  NAND4V2_8TH40 U519 ( .A1(n240), .A2(n241), .A3(n242), .A4(n243), .ZN(
        exe_result_o[9]) );
  AOI221V2_8TH40 U520 ( .A1(cp0_ex_rdata[9]), .A2(n254), .B1(wb_cp0_wdata[9]), 
        .B2(n255), .C(n256), .ZN(n241) );
  AOI221V2_8TH40 U521 ( .A1(N1816), .A2(n262), .B1(n263), .B2(gpr1_data[9]), 
        .C(n264), .ZN(n240) );
  AOI221V2_8TH40 U522 ( .A1(sum_res[9]), .A2(n244), .B1(link_addr[9]), .B2(
        n245), .C(n246), .ZN(n243) );
  NAND4V2_8TH40 U523 ( .A1(n722), .A2(n723), .A3(n724), .A4(n725), .ZN(
        exe_result_o[10]) );
  AOI221V2_8TH40 U524 ( .A1(cp0_ex_rdata[10]), .A2(n254), .B1(wb_cp0_wdata[10]), .B2(n255), .C(n729), .ZN(n723) );
  AOI221V2_8TH40 U525 ( .A1(N1817), .A2(n262), .B1(n263), .B2(gpr1_data[10]), 
        .C(n730), .ZN(n722) );
  AOI221V2_8TH40 U526 ( .A1(sum_res[10]), .A2(n244), .B1(link_addr[10]), .B2(
        n245), .C(n726), .ZN(n725) );
  NAND4V2_8TH40 U527 ( .A1(n712), .A2(n713), .A3(n714), .A4(n715), .ZN(
        exe_result_o[11]) );
  AOI221V2_8TH40 U528 ( .A1(cp0_ex_rdata[11]), .A2(n254), .B1(wb_cp0_wdata[11]), .B2(n255), .C(n718), .ZN(n713) );
  AOI221V2_8TH40 U529 ( .A1(N1818), .A2(n262), .B1(n263), .B2(gpr1_data[11]), 
        .C(n719), .ZN(n712) );
  AOI221V2_8TH40 U530 ( .A1(sum_res[11]), .A2(n244), .B1(link_addr[11]), .B2(
        n245), .C(n716), .ZN(n715) );
  NAND4V2_8TH40 U531 ( .A1(n691), .A2(n692), .A3(n693), .A4(n694), .ZN(
        exe_result_o[13]) );
  AOI221V2_8TH40 U532 ( .A1(cp0_ex_rdata[13]), .A2(n254), .B1(wb_cp0_wdata[13]), .B2(n255), .C(n698), .ZN(n692) );
  AOI221V2_8TH40 U533 ( .A1(N1820), .A2(n262), .B1(n263), .B2(gpr1_data[13]), 
        .C(n699), .ZN(n691) );
  AOI221V2_8TH40 U534 ( .A1(sum_res[13]), .A2(n244), .B1(link_addr[13]), .B2(
        n245), .C(n695), .ZN(n694) );
  NAND4V2_8TH40 U535 ( .A1(n282), .A2(n283), .A3(n284), .A4(n285), .ZN(
        exe_result_o[7]) );
  AOI221V2_8TH40 U536 ( .A1(N1814), .A2(n262), .B1(n263), .B2(gpr1_data[7]), 
        .C(n290), .ZN(n282) );
  AOI222V2_8TH40 U537 ( .A1(wb_cp0_wdata[7]), .A2(n255), .B1(n289), .B2(n1005), 
        .C1(cp0_ex_rdata[7]), .C2(n254), .ZN(n283) );
  AOI222V2_8TH40 U538 ( .A1(n288), .A2(lo[7]), .B1(N1846), .B2(n252), .C1(
        mem_cp0_wdata[7]), .C2(n250), .ZN(n284) );
  NAND4V2_8TH40 U539 ( .A1(n670), .A2(n671), .A3(n672), .A4(n673), .ZN(
        exe_result_o[15]) );
  AOI221V2_8TH40 U540 ( .A1(N1822), .A2(n262), .B1(n263), .B2(gpr1_data[15]), 
        .C(n676), .ZN(n670) );
  AOI222V2_8TH40 U541 ( .A1(wb_cp0_wdata[15]), .A2(n255), .B1(n289), .B2(n997), 
        .C1(cp0_ex_rdata[15]), .C2(n254), .ZN(n671) );
  AOI222V2_8TH40 U542 ( .A1(n288), .A2(lo[15]), .B1(N1854), .B2(n252), .C1(
        mem_cp0_wdata[15]), .C2(n250), .ZN(n672) );
  AOI22V2_8TH40 U543 ( .A1(N1811), .A2(n262), .B1(n263), .B2(gpr1_data[4]), 
        .ZN(n335) );
  NAND4V2_8TH40 U544 ( .A1(n628), .A2(n629), .A3(n630), .A4(n631), .ZN(
        exe_result_o[19]) );
  AOI211V2_8TH40 U545 ( .A1(n263), .A2(gpr1_data[19]), .B(n634), .C(n583), 
        .ZN(n628) );
  AOI222V2_8TH40 U546 ( .A1(N1826), .A2(n262), .B1(cp0_ex_rdata[19]), .B2(n254), .C1(wb_cp0_wdata[19]), .C2(n255), .ZN(n629) );
  NAND4V2_8TH40 U547 ( .A1(n541), .A2(n542), .A3(n543), .A4(n544), .ZN(
        exe_result_o[23]) );
  AOI211V2_8TH40 U548 ( .A1(n263), .A2(gpr1_data[23]), .B(n547), .C(n538), 
        .ZN(n541) );
  AOI222V2_8TH40 U549 ( .A1(N1830), .A2(n262), .B1(cp0_ex_rdata[23]), .B2(n254), .C1(wb_cp0_wdata[23]), .C2(n255), .ZN(n542) );
  NAND4V2_8TH40 U550 ( .A1(n406), .A2(n407), .A3(n408), .A4(n409), .ZN(
        exe_result_o[31]) );
  I2NOR3V2_8TH40 U551 ( .A1(n410), .A2(n411), .B(n412), .ZN(n409) );
  NAND4V2_8TH40 U552 ( .A1(n733), .A2(n734), .A3(n735), .A4(n736), .ZN(
        exe_result_o[0]) );
  I2NOR3V2_8TH40 U553 ( .A1(n737), .A2(n738), .B(n739), .ZN(n736) );
  AOI211V2_8TH40 U554 ( .A1(n326), .A2(n779), .B(n780), .C(n781), .ZN(n735) );
  AOI22V2_8TH40 U555 ( .A1(sum_res[0]), .A2(n244), .B1(link_addr[0]), .B2(n245), .ZN(n734) );
  NAND4V2_8TH40 U556 ( .A1(n236), .A2(inst_type[6]), .A3(n837), .A4(
        inst_type[2]), .ZN(n831) );
  AOI22V2_8TH40 U557 ( .A1(n324), .A2(n612), .B1(sum_res[1]), .B2(n244), .ZN(
        n594) );
  I2NAND4V2_8TH40 U558 ( .A1(n613), .A2(n463), .B1(n614), .B2(n615), .ZN(n612)
         );
  AOI22V2_8TH40 U559 ( .A1(n324), .A2(n456), .B1(sum_res[2]), .B2(n244), .ZN(
        n439) );
  NAND4V2_8TH40 U560 ( .A1(n457), .A2(n458), .A3(n459), .A4(n460), .ZN(n456)
         );
  AOI31V2_8TH40 U561 ( .A1(n464), .A2(n1035), .A3(n465), .B(n466), .ZN(n459)
         );
  NAND4V2_8TH40 U562 ( .A1(n363), .A2(n364), .A3(n365), .A4(n366), .ZN(
        exe_result_o[3]) );
  I2NOR3V2_8TH40 U563 ( .A1(n367), .A2(n368), .B(n369), .ZN(n366) );
  AOI22V2_8TH40 U564 ( .A1(n289), .A2(n1009), .B1(cp0_ex_rdata[3]), .B2(n254), 
        .ZN(n364) );
  AOI22V2_8TH40 U565 ( .A1(wb_cp0_wdata[3]), .A2(n255), .B1(N1810), .B2(n262), 
        .ZN(n363) );
  OAI211V2_8TH40 U566 ( .A1(n912), .A2(n314), .B(n740), .C(n741), .ZN(n739) );
  MUX3V2_8TH40 U567 ( .I0(n316), .I1(n317), .I2(n752), .S0(gpr1_data[0]), .S1(
        gpr2_data[0]), .Z(n740) );
  AOI22V2_8TH40 U568 ( .A1(wb_cp0_wdata[0]), .A2(n255), .B1(N1807), .B2(n262), 
        .ZN(n741) );
  NOR2V2_8TH40 U569 ( .A1(n319), .A2(n753), .ZN(n752) );
  NAND4V2_8TH40 U570 ( .A1(n765), .A2(mem_cp0_we), .A3(n766), .A4(n767), .ZN(
        n750) );
  NOR3V2_8TH40 U571 ( .A1(n768), .A2(n769), .A3(n770), .ZN(n767) );
  AOI22V2_8TH40 U572 ( .A1(n289), .A2(n1012), .B1(cp0_ex_rdata[0]), .B2(n254), 
        .ZN(n737) );
  OAI211V2_8TH40 U573 ( .A1(n1021), .A2(n314), .B(n476), .C(n523), .ZN(n522)
         );
  MUX3V2_8TH40 U574 ( .I0(n316), .I1(n317), .I2(n524), .S0(gpr1_data[25]), 
        .S1(gpr2_data[25]), .Z(n523) );
  NOR2V2_8TH40 U575 ( .A1(n319), .A2(n525), .ZN(n524) );
  OAI211V2_8TH40 U576 ( .A1(n1026), .A2(n314), .B(n558), .C(n580), .ZN(n579)
         );
  MUX3V2_8TH40 U577 ( .I0(n316), .I1(n317), .I2(n581), .S0(gpr1_data[20]), 
        .S1(gpr2_data[20]), .Z(n580) );
  NOR2V2_8TH40 U578 ( .A1(n319), .A2(n582), .ZN(n581) );
  OAI211V2_8TH40 U579 ( .A1(n1024), .A2(n314), .B(n558), .C(n559), .ZN(n557)
         );
  MUX3V2_8TH40 U580 ( .I0(n316), .I1(n317), .I2(n560), .S0(gpr1_data[22]), 
        .S1(gpr2_data[22]), .Z(n559) );
  NOR2V2_8TH40 U581 ( .A1(n319), .A2(n561), .ZN(n560) );
  OAI211V2_8TH40 U582 ( .A1(n1020), .A2(n314), .B(n476), .C(n512), .ZN(n511)
         );
  MUX3V2_8TH40 U583 ( .I0(n316), .I1(n317), .I2(n513), .S0(gpr1_data[26]), 
        .S1(gpr2_data[26]), .Z(n512) );
  NOR2V2_8TH40 U584 ( .A1(n319), .A2(n514), .ZN(n513) );
  OAI211V2_8TH40 U585 ( .A1(n1019), .A2(n314), .B(n476), .C(n500), .ZN(n499)
         );
  MUX3V2_8TH40 U586 ( .I0(n316), .I1(n317), .I2(n501), .S0(gpr1_data[27]), 
        .S1(gpr2_data[27]), .Z(n500) );
  NOR2V2_8TH40 U587 ( .A1(n319), .A2(n502), .ZN(n501) );
  OAI211V2_8TH40 U588 ( .A1(n1022), .A2(n314), .B(n476), .C(n535), .ZN(n534)
         );
  MUX3V2_8TH40 U589 ( .I0(n316), .I1(n317), .I2(n536), .S0(gpr1_data[24]), 
        .S1(gpr2_data[24]), .Z(n535) );
  NOR2V2_8TH40 U590 ( .A1(n319), .A2(n537), .ZN(n536) );
  OAI211V2_8TH40 U591 ( .A1(n1017), .A2(n314), .B(n476), .C(n477), .ZN(n475)
         );
  MUX3V2_8TH40 U592 ( .I0(n316), .I1(n317), .I2(n478), .S0(gpr1_data[29]), 
        .S1(gpr2_data[29]), .Z(n477) );
  NOR2V2_8TH40 U593 ( .A1(n319), .A2(n479), .ZN(n478) );
  OAI211V2_8TH40 U594 ( .A1(n370), .A2(n346), .B(n371), .C(n372), .ZN(n369) );
  OAI31V2_8TH40 U595 ( .A1(n373), .A2(n374), .A3(n375), .B(n326), .ZN(n371) );
  AOI211V2_8TH40 U596 ( .A1(n383), .A2(n1023), .B(n384), .C(n385), .ZN(n370)
         );
  AOI22V2_8TH40 U597 ( .A1(sum_res[3]), .A2(n244), .B1(link_addr[3]), .B2(n245), .ZN(n372) );
  INOR2V2_8TH40 U598 ( .A1(n828), .B1(n829), .ZN(except_type_o[11]) );
  NAND4V2_8TH40 U599 ( .A1(n771), .A2(wb_cp0_we), .A3(n772), .A4(n773), .ZN(
        n751) );
  NOR3V2_8TH40 U600 ( .A1(n774), .A2(n775), .A3(n776), .ZN(n773) );
  AOI22V2_8TH40 U601 ( .A1(n328), .A2(n526), .B1(n326), .B2(n596), .ZN(n595)
         );
  NAND4V2_8TH40 U602 ( .A1(n597), .A2(n598), .A3(n599), .A4(n600), .ZN(n596)
         );
  AOI211V2_8TH40 U603 ( .A1(n601), .A2(gpr1_data[12]), .B(n602), .C(n449), 
        .ZN(n600) );
  AOI22V2_8TH40 U604 ( .A1(n441), .A2(n328), .B1(n326), .B2(n442), .ZN(n440)
         );
  NAND4V2_8TH40 U605 ( .A1(n443), .A2(n400), .A3(n444), .A4(n445), .ZN(n442)
         );
  AOI33V2_8TH40 U606 ( .A1(gpr1_data[19]), .A2(n1026), .A3(n450), .B1(n451), 
        .B2(n452), .B3(n453), .ZN(n444) );
  AOI31V2_8TH40 U607 ( .A1(n782), .A2(n390), .A3(n783), .B(n346), .ZN(n781) );
  AOI211V2_8TH40 U608 ( .A1(n785), .A2(n625), .B(n397), .C(n617), .ZN(n783) );
  OAI21V2_8TH40 U609 ( .A1(n1041), .A2(n314), .B(n315), .ZN(n313) );
  MUX3V2_8TH40 U610 ( .I0(n316), .I1(n317), .I2(n318), .S0(gpr1_data[5]), .S1(
        gpr2_data[5]), .Z(n315) );
  NOR2V2_8TH40 U611 ( .A1(n319), .A2(n320), .ZN(n318) );
  OAI21V2_8TH40 U612 ( .A1(n353), .A2(n299), .B(n354), .ZN(n342) );
  AO31V2_8TH40 U613 ( .A1(n355), .A2(n356), .A3(n357), .B(n358), .Z(n354) );
  NAND4V2_8TH40 U614 ( .A1(n597), .A2(n400), .A3(n795), .A4(n796), .ZN(n779)
         );
  AOAOAOI211111V2_8TH40 U615 ( .A1(gpr1_data[26]), .A2(n1019), .B(
        gpr1_data[28]), .C(n1017), .D(gpr1_data[30]), .E(n1015), .F(n799), 
        .ZN(n795) );
  AOI21V2_8TH40 U616 ( .A1(n344), .A2(n345), .B(n346), .ZN(n343) );
  AOI32V2_8TH40 U617 ( .A1(gpr1_data[16]), .A2(n1031), .A3(n347), .B1(n348), 
        .B2(n349), .ZN(n345) );
  NOR2V2_8TH40 U618 ( .A1(n319), .A2(n591), .ZN(n590) );
  NOR2V2_8TH40 U619 ( .A1(n319), .A2(n436), .ZN(n435) );
  NAND3V2_8TH40 U620 ( .A1(n788), .A2(n789), .A3(n389), .ZN(n352) );
  AO211V2_8TH40 U621 ( .A1(gpr1_data[14]), .A2(n360), .B(n797), .C(n798), .Z(
        n361) );
  MUX3V2_8TH40 U622 ( .I0(n265), .I1(n266), .I2(n709), .S0(gpr1_data[12]), 
        .S1(gpr2_data[12]), .Z(n708) );
  NAND2V2_8TH40 U623 ( .A1(n710), .A2(n269), .ZN(n709) );
  MUX3V2_8TH40 U624 ( .I0(n265), .I1(n266), .I2(n686), .S0(gpr1_data[14]), 
        .S1(gpr2_data[14]), .Z(n685) );
  NAND2V2_8TH40 U625 ( .A1(n687), .A2(n269), .ZN(n686) );
  MUX3V2_8TH40 U626 ( .I0(n265), .I1(n266), .I2(n339), .S0(gpr1_data[4]), .S1(
        gpr2_data[4]), .Z(n338) );
  NAND2V2_8TH40 U627 ( .A1(n340), .A2(n269), .ZN(n339) );
  MUX3V2_8TH40 U628 ( .I0(n265), .I1(n266), .I2(n636), .S0(gpr1_data[19]), 
        .S1(gpr2_data[19]), .Z(n634) );
  NAND2V2_8TH40 U629 ( .A1(n637), .A2(n269), .ZN(n636) );
  MUX3V2_8TH40 U630 ( .I0(n265), .I1(n266), .I2(n549), .S0(gpr1_data[23]), 
        .S1(gpr2_data[23]), .Z(n547) );
  NAND2V2_8TH40 U631 ( .A1(n550), .A2(n269), .ZN(n549) );
  MUX3V2_8TH40 U632 ( .I0(n265), .I1(n266), .I2(n304), .S0(gpr1_data[6]), .S1(
        gpr2_data[6]), .Z(n303) );
  NAND2V2_8TH40 U633 ( .A1(n305), .A2(n269), .ZN(n304) );
  MUX3V2_8TH40 U634 ( .I0(n265), .I1(n266), .I2(n291), .S0(gpr1_data[7]), .S1(
        gpr2_data[7]), .Z(n290) );
  NAND2V2_8TH40 U635 ( .A1(n292), .A2(n269), .ZN(n291) );
  MUX3V2_8TH40 U636 ( .I0(n265), .I1(n266), .I2(n280), .S0(gpr1_data[8]), .S1(
        gpr2_data[8]), .Z(n279) );
  NAND2V2_8TH40 U637 ( .A1(n281), .A2(n269), .ZN(n280) );
  MUX3V2_8TH40 U638 ( .I0(n265), .I1(n266), .I2(n267), .S0(gpr1_data[9]), .S1(
        gpr2_data[9]), .Z(n264) );
  NAND2V2_8TH40 U639 ( .A1(n268), .A2(n269), .ZN(n267) );
  MUX3V2_8TH40 U640 ( .I0(n265), .I1(n266), .I2(n731), .S0(gpr1_data[10]), 
        .S1(gpr2_data[10]), .Z(n730) );
  NAND2V2_8TH40 U641 ( .A1(n732), .A2(n269), .ZN(n731) );
  MUX3V2_8TH40 U642 ( .I0(n265), .I1(n266), .I2(n720), .S0(gpr1_data[11]), 
        .S1(gpr2_data[11]), .Z(n719) );
  NAND2V2_8TH40 U643 ( .A1(n721), .A2(n269), .ZN(n720) );
  MUX3V2_8TH40 U644 ( .I0(n265), .I1(n266), .I2(n700), .S0(gpr1_data[13]), 
        .S1(gpr2_data[13]), .Z(n699) );
  NAND2V2_8TH40 U645 ( .A1(n701), .A2(n269), .ZN(n700) );
  MUX3V2_8TH40 U646 ( .I0(n265), .I1(n266), .I2(n677), .S0(gpr1_data[15]), 
        .S1(gpr2_data[15]), .Z(n676) );
  NAND2V2_8TH40 U647 ( .A1(n678), .A2(n269), .ZN(n677) );
  MUX3V2_8TH40 U648 ( .I0(n265), .I1(n266), .I2(n668), .S0(gpr1_data[16]), 
        .S1(gpr2_data[16]), .Z(n667) );
  NAND2V2_8TH40 U649 ( .A1(n669), .A2(n269), .ZN(n668) );
  MUX3V2_8TH40 U650 ( .I0(n265), .I1(n266), .I2(n657), .S0(gpr1_data[17]), 
        .S1(gpr2_data[17]), .Z(n656) );
  NAND2V2_8TH40 U651 ( .A1(n658), .A2(n269), .ZN(n657) );
  MUX3V2_8TH40 U652 ( .I0(n265), .I1(n266), .I2(n647), .S0(gpr1_data[18]), 
        .S1(gpr2_data[18]), .Z(n646) );
  NAND2V2_8TH40 U653 ( .A1(n648), .A2(n269), .ZN(n647) );
  MUX3V2_8TH40 U654 ( .I0(n265), .I1(n266), .I2(n571), .S0(gpr1_data[21]), 
        .S1(gpr2_data[21]), .Z(n570) );
  NAND2V2_8TH40 U655 ( .A1(n572), .A2(n269), .ZN(n571) );
  MUX3V2_8TH40 U656 ( .I0(n265), .I1(n266), .I2(n491), .S0(gpr1_data[28]), 
        .S1(gpr2_data[28]), .Z(n490) );
  NAND2V2_8TH40 U657 ( .A1(n492), .A2(n269), .ZN(n491) );
  MUX3V2_8TH40 U658 ( .I0(n265), .I1(n266), .I2(n428), .S0(gpr1_data[30]), 
        .S1(gpr2_data[30]), .Z(n427) );
  NAND2V2_8TH40 U659 ( .A1(n429), .A2(n269), .ZN(n428) );
  NOR2V0_8TH40 U660 ( .A1(n3), .A2(n41), .ZN(n121) );
  OAI211V2_8TH40 U661 ( .A1(n21), .A2(n37), .B(n187), .C(n188), .ZN(hi_o[21])
         );
  OAI211V2_8TH40 U662 ( .A1(n183), .A2(n37), .B(n184), .C(n185), .ZN(hi_o[22])
         );
  OAI211V2_8TH40 U663 ( .A1(n179), .A2(n37), .B(n180), .C(n181), .ZN(hi_o[23])
         );
  OAI211V2_8TH40 U664 ( .A1(n175), .A2(n37), .B(n176), .C(n177), .ZN(hi_o[24])
         );
  OAI211V2_8TH40 U665 ( .A1(n171), .A2(n37), .B(n172), .C(n173), .ZN(hi_o[25])
         );
  OAI211V2_8TH40 U666 ( .A1(n167), .A2(n37), .B(n168), .C(n169), .ZN(hi_o[26])
         );
  OAI211V2_8TH40 U667 ( .A1(n163), .A2(n37), .B(n164), .C(n165), .ZN(hi_o[27])
         );
  OAI211V2_8TH40 U668 ( .A1(n20), .A2(n37), .B(n160), .C(n161), .ZN(hi_o[28])
         );
  OAI211V2_8TH40 U669 ( .A1(n156), .A2(n37), .B(n157), .C(n158), .ZN(hi_o[29])
         );
  OAI211V2_8TH40 U670 ( .A1(n19), .A2(n37), .B(n150), .C(n151), .ZN(hi_o[30])
         );
  OAI211V2_8TH40 U671 ( .A1(n146), .A2(n37), .B(n147), .C(n148), .ZN(hi_o[31])
         );
  OAI33V2_8TH40 U672 ( .A1(n812), .A2(inst_type[4]), .A3(n813), .B1(n814), 
        .B2(n815), .B3(n816), .ZN(except_type_o[10]) );
  AOAI211V2_8TH40 U673 ( .A1(n817), .A2(n810), .B(n818), .C(n777), .ZN(n814)
         );
  AND2V2_8TH40 U674 ( .A1(n912), .A2(n913), .Z(n4) );
  AND2V2_8TH40 U675 ( .A1(n4), .A2(n914), .Z(n15) );
  AND2V2_8TH40 U676 ( .A1(n15), .A2(n915), .Z(n16) );
  AND2V2_8TH40 U677 ( .A1(n16), .A2(n916), .Z(n17) );
  XOR2V2_8TH40 U678 ( .A1(n912), .A2(n913), .Z(N1872) );
  XOR2V2_8TH40 U679 ( .A1(n4), .A2(n914), .Z(N1873) );
  XOR2V2_8TH40 U680 ( .A1(n16), .A2(n916), .Z(N1875) );
  NOR2V0P5_8TH40 U681 ( .A1(inst_type[0]), .A2(n18), .ZN(signed_div) );
  CLKNV1_8TH40 U682 ( .I(n19), .ZN(n982) );
  CLKNV1_8TH40 U683 ( .I(n20), .ZN(n984) );
  CLKNV1_8TH40 U684 ( .I(n21), .ZN(n991) );
  CLKNV1_8TH40 U685 ( .I(n22), .ZN(n994) );
  CLKNV1_8TH40 U686 ( .I(n23), .ZN(n995) );
  CLKNV1_8TH40 U687 ( .I(n24), .ZN(n996) );
  CLKNV1_8TH40 U688 ( .I(n25), .ZN(n999) );
  CLKNV1_8TH40 U689 ( .I(n26), .ZN(n1001) );
  CLKNV1_8TH40 U690 ( .I(n27), .ZN(n1002) );
  CLKNV1_8TH40 U691 ( .I(n28), .ZN(n1003) );
  CLKNV1_8TH40 U692 ( .I(n29), .ZN(n1004) );
  CLKNV1_8TH40 U693 ( .I(n30), .ZN(n1006) );
  CLKNV1_8TH40 U694 ( .I(n31), .ZN(n1008) );
  CLKNV1_8TH40 U695 ( .I(n32), .ZN(n1010) );
  CLKNV1_8TH40 U696 ( .I(n33), .ZN(n1011) );
  CKMUX2V2_8TH40 U697 ( .I0(gpr2_data[9]), .I1(N574), .S(n34), .Z(
        mul_opdata2[9]) );
  CKMUX2V2_8TH40 U698 ( .I0(gpr2_data[8]), .I1(N573), .S(n34), .Z(
        mul_opdata2[8]) );
  CKMUX2V2_8TH40 U699 ( .I0(gpr2_data[7]), .I1(N572), .S(n34), .Z(
        mul_opdata2[7]) );
  CKMUX2V2_8TH40 U700 ( .I0(gpr2_data[6]), .I1(N571), .S(n34), .Z(
        mul_opdata2[6]) );
  CKMUX2V2_8TH40 U701 ( .I0(gpr2_data[5]), .I1(N570), .S(n34), .Z(
        mul_opdata2[5]) );
  CKMUX2V2_8TH40 U702 ( .I0(gpr2_data[4]), .I1(N569), .S(n34), .Z(
        mul_opdata2[4]) );
  CKMUX2V2_8TH40 U703 ( .I0(gpr2_data[3]), .I1(N568), .S(n34), .Z(
        mul_opdata2[3]) );
  CKMUX2V2_8TH40 U704 ( .I0(gpr2_data[31]), .I1(N596), .S(n34), .Z(
        mul_opdata2[31]) );
  CKMUX2V2_8TH40 U705 ( .I0(gpr2_data[30]), .I1(N595), .S(n34), .Z(
        mul_opdata2[30]) );
  CKMUX2V2_8TH40 U706 ( .I0(gpr2_data[2]), .I1(N567), .S(n34), .Z(
        mul_opdata2[2]) );
  CKMUX2V2_8TH40 U707 ( .I0(gpr2_data[29]), .I1(N594), .S(n34), .Z(
        mul_opdata2[29]) );
  CKMUX2V2_8TH40 U708 ( .I0(gpr2_data[28]), .I1(N593), .S(n34), .Z(
        mul_opdata2[28]) );
  CKMUX2V2_8TH40 U709 ( .I0(gpr2_data[27]), .I1(N592), .S(n34), .Z(
        mul_opdata2[27]) );
  CKMUX2V2_8TH40 U710 ( .I0(gpr2_data[26]), .I1(N591), .S(n34), .Z(
        mul_opdata2[26]) );
  CKMUX2V2_8TH40 U711 ( .I0(gpr2_data[25]), .I1(N590), .S(n34), .Z(
        mul_opdata2[25]) );
  CKMUX2V2_8TH40 U712 ( .I0(gpr2_data[24]), .I1(N589), .S(n34), .Z(
        mul_opdata2[24]) );
  CKMUX2V2_8TH40 U713 ( .I0(gpr2_data[23]), .I1(N588), .S(n34), .Z(
        mul_opdata2[23]) );
  CKMUX2V2_8TH40 U714 ( .I0(gpr2_data[22]), .I1(N587), .S(n34), .Z(
        mul_opdata2[22]) );
  CKMUX2V2_8TH40 U715 ( .I0(gpr2_data[21]), .I1(N586), .S(n34), .Z(
        mul_opdata2[21]) );
  CKMUX2V2_8TH40 U716 ( .I0(gpr2_data[20]), .I1(N585), .S(n34), .Z(
        mul_opdata2[20]) );
  CKMUX2V2_8TH40 U717 ( .I0(gpr2_data[1]), .I1(N566), .S(n34), .Z(
        mul_opdata2[1]) );
  CKMUX2V2_8TH40 U718 ( .I0(gpr2_data[19]), .I1(N584), .S(n34), .Z(
        mul_opdata2[19]) );
  CKMUX2V2_8TH40 U719 ( .I0(gpr2_data[18]), .I1(N583), .S(n34), .Z(
        mul_opdata2[18]) );
  CKMUX2V2_8TH40 U720 ( .I0(gpr2_data[17]), .I1(N582), .S(n34), .Z(
        mul_opdata2[17]) );
  CKMUX2V2_8TH40 U721 ( .I0(gpr2_data[16]), .I1(N581), .S(n34), .Z(
        mul_opdata2[16]) );
  CKMUX2V2_8TH40 U722 ( .I0(gpr2_data[15]), .I1(N580), .S(n34), .Z(
        mul_opdata2[15]) );
  CKMUX2V2_8TH40 U723 ( .I0(gpr2_data[14]), .I1(N579), .S(n34), .Z(
        mul_opdata2[14]) );
  CKMUX2V2_8TH40 U724 ( .I0(gpr2_data[13]), .I1(N578), .S(n34), .Z(
        mul_opdata2[13]) );
  CKMUX2V2_8TH40 U725 ( .I0(gpr2_data[12]), .I1(N577), .S(n34), .Z(
        mul_opdata2[12]) );
  CKMUX2V2_8TH40 U726 ( .I0(gpr2_data[11]), .I1(N576), .S(n34), .Z(
        mul_opdata2[11]) );
  CKMUX2V2_8TH40 U727 ( .I0(gpr2_data[10]), .I1(N575), .S(n34), .Z(
        mul_opdata2[10]) );
  CKMUX2V2_8TH40 U728 ( .I0(gpr2_data[0]), .I1(N565), .S(n34), .Z(
        mul_opdata2[0]) );
  CKMUX2V2_8TH40 U729 ( .I0(gpr1_data[9]), .I1(N509), .S(n36), .Z(
        mul_opdata1[9]) );
  CKMUX2V2_8TH40 U730 ( .I0(gpr1_data[8]), .I1(N508), .S(n36), .Z(
        mul_opdata1[8]) );
  CKMUX2V2_8TH40 U731 ( .I0(gpr1_data[7]), .I1(N507), .S(n36), .Z(
        mul_opdata1[7]) );
  CKMUX2V2_8TH40 U732 ( .I0(gpr1_data[6]), .I1(N506), .S(n36), .Z(
        mul_opdata1[6]) );
  CKMUX2V2_8TH40 U733 ( .I0(gpr1_data[5]), .I1(N505), .S(n36), .Z(
        mul_opdata1[5]) );
  CKMUX2V2_8TH40 U734 ( .I0(gpr1_data[4]), .I1(N504), .S(n36), .Z(
        mul_opdata1[4]) );
  CKMUX2V2_8TH40 U735 ( .I0(gpr1_data[3]), .I1(N503), .S(n36), .Z(
        mul_opdata1[3]) );
  CKMUX2V2_8TH40 U736 ( .I0(gpr1_data[31]), .I1(N531), .S(n36), .Z(
        mul_opdata1[31]) );
  CKMUX2V2_8TH40 U737 ( .I0(gpr1_data[30]), .I1(N530), .S(n36), .Z(
        mul_opdata1[30]) );
  CKMUX2V2_8TH40 U738 ( .I0(gpr1_data[2]), .I1(N502), .S(n36), .Z(
        mul_opdata1[2]) );
  CKMUX2V2_8TH40 U739 ( .I0(gpr1_data[29]), .I1(N529), .S(n36), .Z(
        mul_opdata1[29]) );
  CKMUX2V2_8TH40 U740 ( .I0(gpr1_data[28]), .I1(N528), .S(n36), .Z(
        mul_opdata1[28]) );
  CKMUX2V2_8TH40 U741 ( .I0(gpr1_data[27]), .I1(N527), .S(n36), .Z(
        mul_opdata1[27]) );
  CKMUX2V2_8TH40 U742 ( .I0(gpr1_data[26]), .I1(N526), .S(n36), .Z(
        mul_opdata1[26]) );
  CKMUX2V2_8TH40 U743 ( .I0(gpr1_data[25]), .I1(N525), .S(n36), .Z(
        mul_opdata1[25]) );
  CKMUX2V2_8TH40 U744 ( .I0(gpr1_data[24]), .I1(N524), .S(n36), .Z(
        mul_opdata1[24]) );
  CKMUX2V2_8TH40 U745 ( .I0(gpr1_data[23]), .I1(N523), .S(n36), .Z(
        mul_opdata1[23]) );
  CKMUX2V2_8TH40 U746 ( .I0(gpr1_data[22]), .I1(N522), .S(n36), .Z(
        mul_opdata1[22]) );
  CKMUX2V2_8TH40 U747 ( .I0(gpr1_data[21]), .I1(N521), .S(n36), .Z(
        mul_opdata1[21]) );
  CKMUX2V2_8TH40 U748 ( .I0(gpr1_data[20]), .I1(N520), .S(n36), .Z(
        mul_opdata1[20]) );
  CKMUX2V2_8TH40 U749 ( .I0(gpr1_data[1]), .I1(N501), .S(n36), .Z(
        mul_opdata1[1]) );
  CKMUX2V2_8TH40 U750 ( .I0(gpr1_data[19]), .I1(N519), .S(n36), .Z(
        mul_opdata1[19]) );
  CKMUX2V2_8TH40 U751 ( .I0(gpr1_data[18]), .I1(N518), .S(n36), .Z(
        mul_opdata1[18]) );
  CKMUX2V2_8TH40 U752 ( .I0(gpr1_data[17]), .I1(N517), .S(n36), .Z(
        mul_opdata1[17]) );
  CKMUX2V2_8TH40 U753 ( .I0(gpr1_data[16]), .I1(N516), .S(n36), .Z(
        mul_opdata1[16]) );
  CKMUX2V2_8TH40 U754 ( .I0(gpr1_data[15]), .I1(N515), .S(n36), .Z(
        mul_opdata1[15]) );
  CKMUX2V2_8TH40 U755 ( .I0(gpr1_data[14]), .I1(N514), .S(n36), .Z(
        mul_opdata1[14]) );
  CKMUX2V2_8TH40 U756 ( .I0(gpr1_data[13]), .I1(N513), .S(n36), .Z(
        mul_opdata1[13]) );
  CKMUX2V2_8TH40 U757 ( .I0(gpr1_data[12]), .I1(N512), .S(n36), .Z(
        mul_opdata1[12]) );
  CKMUX2V2_8TH40 U758 ( .I0(gpr1_data[11]), .I1(N511), .S(n36), .Z(
        mul_opdata1[11]) );
  CKMUX2V2_8TH40 U759 ( .I0(gpr1_data[10]), .I1(N510), .S(n36), .Z(
        mul_opdata1[10]) );
  CKMUX2V2_8TH40 U760 ( .I0(gpr1_data[0]), .I1(N500), .S(n36), .Z(
        mul_opdata1[0]) );
  AOI22V0_8TH40 U761 ( .A1(n41), .A2(n972), .B1(n42), .B2(lo[9]), .ZN(n38) );
  AOI22V0_8TH40 U762 ( .A1(n41), .A2(n973), .B1(n42), .B2(lo[8]), .ZN(n43) );
  AOI22V0_8TH40 U763 ( .A1(n41), .A2(n974), .B1(n42), .B2(lo[7]), .ZN(n45) );
  AOI22V0_8TH40 U764 ( .A1(n41), .A2(n975), .B1(n42), .B2(lo[6]), .ZN(n47) );
  AOI22V0_8TH40 U765 ( .A1(n41), .A2(n976), .B1(n42), .B2(lo[5]), .ZN(n49) );
  AOI22V0_8TH40 U766 ( .A1(n41), .A2(n977), .B1(n42), .B2(lo[4]), .ZN(n51) );
  AOI22V0_8TH40 U767 ( .A1(n41), .A2(n978), .B1(n42), .B2(lo[3]), .ZN(n53) );
  AOI22V0_8TH40 U768 ( .A1(n41), .A2(n950), .B1(n42), .B2(lo[31]), .ZN(n55) );
  AOI22V0_8TH40 U769 ( .A1(n41), .A2(n951), .B1(n42), .B2(lo[30]), .ZN(n57) );
  AOI22V0_8TH40 U770 ( .A1(n41), .A2(n979), .B1(n42), .B2(lo[2]), .ZN(n59) );
  AOI22V0_8TH40 U771 ( .A1(n41), .A2(n952), .B1(n42), .B2(lo[29]), .ZN(n61) );
  AOI22V0_8TH40 U772 ( .A1(n41), .A2(n953), .B1(n42), .B2(lo[28]), .ZN(n63) );
  AOI22V0_8TH40 U773 ( .A1(n41), .A2(n954), .B1(n42), .B2(lo[27]), .ZN(n65) );
  AOI22V0_8TH40 U774 ( .A1(n41), .A2(n955), .B1(n42), .B2(lo[26]), .ZN(n67) );
  AOI22V0_8TH40 U775 ( .A1(n41), .A2(n956), .B1(n42), .B2(lo[25]), .ZN(n69) );
  AOI22V0_8TH40 U776 ( .A1(n41), .A2(n957), .B1(n42), .B2(lo[24]), .ZN(n71) );
  AOI22V0_8TH40 U777 ( .A1(n41), .A2(n958), .B1(n42), .B2(lo[23]), .ZN(n73) );
  AOI22V0_8TH40 U778 ( .A1(n41), .A2(n959), .B1(n42), .B2(lo[22]), .ZN(n75) );
  AOI22V0_8TH40 U779 ( .A1(n41), .A2(n960), .B1(n42), .B2(lo[21]), .ZN(n77) );
  AOI22V0_8TH40 U780 ( .A1(n41), .A2(n961), .B1(n42), .B2(lo[20]), .ZN(n79) );
  AOI22V0_8TH40 U781 ( .A1(n41), .A2(n980), .B1(n42), .B2(lo[1]), .ZN(n81) );
  AOI22V0_8TH40 U782 ( .A1(n41), .A2(n962), .B1(n42), .B2(lo[19]), .ZN(n83) );
  AOI22V0_8TH40 U783 ( .A1(n41), .A2(n963), .B1(n42), .B2(lo[18]), .ZN(n85) );
  AOI22V0_8TH40 U784 ( .A1(n41), .A2(n964), .B1(n42), .B2(lo[17]), .ZN(n87) );
  AOI22V0_8TH40 U785 ( .A1(n41), .A2(n965), .B1(n42), .B2(lo[16]), .ZN(n89) );
  AOI22V0_8TH40 U786 ( .A1(n41), .A2(n966), .B1(n42), .B2(lo[15]), .ZN(n91) );
  AOI22V0_8TH40 U787 ( .A1(n41), .A2(n967), .B1(n42), .B2(lo[14]), .ZN(n93) );
  AOI22V0_8TH40 U788 ( .A1(n41), .A2(n968), .B1(n42), .B2(lo[13]), .ZN(n95) );
  AOI22V0_8TH40 U789 ( .A1(n41), .A2(n969), .B1(n42), .B2(lo[12]), .ZN(n97) );
  AOI22V0_8TH40 U790 ( .A1(n41), .A2(n970), .B1(n42), .B2(lo[11]), .ZN(n99) );
  AOI22V0_8TH40 U791 ( .A1(n41), .A2(n971), .B1(n42), .B2(lo[10]), .ZN(n101)
         );
  AOI22V0_8TH40 U792 ( .A1(n41), .A2(n1013), .B1(n42), .B2(lo[0]), .ZN(n103)
         );
  CLKNV1_8TH40 U793 ( .I(n105), .ZN(lo[9]) );
  CLKNV1_8TH40 U794 ( .I(n106), .ZN(lo[8]) );
  CLKNV1_8TH40 U795 ( .I(n107), .ZN(lo[6]) );
  CLKNV1_8TH40 U796 ( .I(n108), .ZN(lo[4]) );
  CLKNV1_8TH40 U797 ( .I(n109), .ZN(lo[30]) );
  CLKNV1_8TH40 U798 ( .I(n110), .ZN(lo[2]) );
  CLKNV1_8TH40 U799 ( .I(n111), .ZN(lo[28]) );
  CLKNV1_8TH40 U800 ( .I(n112), .ZN(lo[21]) );
  CLKNV1_8TH40 U801 ( .I(n113), .ZN(lo[1]) );
  CLKNV1_8TH40 U802 ( .I(n114), .ZN(lo[18]) );
  CLKNV1_8TH40 U803 ( .I(n115), .ZN(lo[17]) );
  CLKNV1_8TH40 U804 ( .I(n116), .ZN(lo[16]) );
  CLKNV1_8TH40 U805 ( .I(n117), .ZN(lo[13]) );
  CLKNV1_8TH40 U806 ( .I(n118), .ZN(lo[11]) );
  CLKNV1_8TH40 U807 ( .I(n119), .ZN(lo[10]) );
  AOI22V0_8TH40 U808 ( .A1(n41), .A2(n940), .B1(n42), .B2(gpr1_data[9]), .ZN(
        n122) );
  CLKNV1_8TH40 U809 ( .I(n124), .ZN(n940) );
  AOI22V0_8TH40 U810 ( .A1(n41), .A2(n941), .B1(n42), .B2(gpr1_data[8]), .ZN(
        n125) );
  CLKNV1_8TH40 U811 ( .I(n127), .ZN(n941) );
  AOI22V0_8TH40 U812 ( .A1(n41), .A2(n942), .B1(n42), .B2(gpr1_data[7]), .ZN(
        n129) );
  CLKNV1_8TH40 U813 ( .I(n131), .ZN(n942) );
  AOI22V0_8TH40 U814 ( .A1(n41), .A2(n943), .B1(n42), .B2(gpr1_data[6]), .ZN(
        n132) );
  CLKNV1_8TH40 U815 ( .I(n134), .ZN(n943) );
  AOI22V0_8TH40 U816 ( .A1(n41), .A2(n944), .B1(n42), .B2(gpr1_data[5]), .ZN(
        n136) );
  CLKNV1_8TH40 U817 ( .I(n138), .ZN(n944) );
  AOI22V0_8TH40 U818 ( .A1(n41), .A2(n945), .B1(n42), .B2(gpr1_data[4]), .ZN(
        n139) );
  CLKNV1_8TH40 U819 ( .I(n141), .ZN(n945) );
  AOI22V0_8TH40 U820 ( .A1(n41), .A2(n946), .B1(n42), .B2(gpr1_data[3]), .ZN(
        n143) );
  CLKNV1_8TH40 U821 ( .I(n145), .ZN(n946) );
  AOI22V0_8TH40 U822 ( .A1(div_res[63]), .A2(n40), .B1(mul_res_tmp1[63]), .B2(
        n3), .ZN(n148) );
  AOI22V0_8TH40 U823 ( .A1(n41), .A2(n918), .B1(n42), .B2(gpr1_data[31]), .ZN(
        n147) );
  CLKNV1_8TH40 U824 ( .I(n149), .ZN(n918) );
  AOI22V0_8TH40 U825 ( .A1(div_res[62]), .A2(n40), .B1(mul_res_tmp1[62]), .B2(
        n3), .ZN(n151) );
  AOI22V0_8TH40 U826 ( .A1(n41), .A2(n919), .B1(n42), .B2(gpr1_data[30]), .ZN(
        n150) );
  CLKNV1_8TH40 U827 ( .I(n152), .ZN(n919) );
  AOI22V0_8TH40 U828 ( .A1(n41), .A2(n947), .B1(n42), .B2(gpr1_data[2]), .ZN(
        n153) );
  CLKNV1_8TH40 U829 ( .I(n155), .ZN(n947) );
  AOI22V0_8TH40 U830 ( .A1(div_res[61]), .A2(n40), .B1(mul_res_tmp1[61]), .B2(
        n3), .ZN(n158) );
  AOI22V0_8TH40 U831 ( .A1(n41), .A2(n920), .B1(n42), .B2(gpr1_data[29]), .ZN(
        n157) );
  CLKNV1_8TH40 U832 ( .I(n159), .ZN(n920) );
  AOI22V0_8TH40 U833 ( .A1(div_res[60]), .A2(n40), .B1(mul_res_tmp1[60]), .B2(
        n3), .ZN(n161) );
  AOI22V0_8TH40 U834 ( .A1(n41), .A2(n921), .B1(n42), .B2(gpr1_data[28]), .ZN(
        n160) );
  CLKNV1_8TH40 U835 ( .I(n162), .ZN(n921) );
  AOI22V0_8TH40 U836 ( .A1(div_res[59]), .A2(n40), .B1(mul_res_tmp1[59]), .B2(
        n3), .ZN(n165) );
  AOI22V0_8TH40 U837 ( .A1(n41), .A2(n922), .B1(n42), .B2(gpr1_data[27]), .ZN(
        n164) );
  CLKNV1_8TH40 U838 ( .I(n166), .ZN(n922) );
  AOI22V0_8TH40 U839 ( .A1(div_res[58]), .A2(n40), .B1(mul_res_tmp1[58]), .B2(
        n3), .ZN(n169) );
  AOI22V0_8TH40 U840 ( .A1(n41), .A2(n923), .B1(n42), .B2(gpr1_data[26]), .ZN(
        n168) );
  CLKNV1_8TH40 U841 ( .I(n170), .ZN(n923) );
  AOI22V0_8TH40 U842 ( .A1(div_res[57]), .A2(n40), .B1(mul_res_tmp1[57]), .B2(
        n3), .ZN(n173) );
  AOI22V0_8TH40 U843 ( .A1(n41), .A2(n924), .B1(n42), .B2(gpr1_data[25]), .ZN(
        n172) );
  CLKNV1_8TH40 U844 ( .I(n174), .ZN(n924) );
  AOI22V0_8TH40 U845 ( .A1(div_res[56]), .A2(n40), .B1(mul_res_tmp1[56]), .B2(
        n3), .ZN(n177) );
  AOI22V0_8TH40 U846 ( .A1(n41), .A2(n925), .B1(n42), .B2(gpr1_data[24]), .ZN(
        n176) );
  CLKNV1_8TH40 U847 ( .I(n178), .ZN(n925) );
  AOI22V0_8TH40 U848 ( .A1(div_res[55]), .A2(n40), .B1(mul_res_tmp1[55]), .B2(
        n3), .ZN(n181) );
  AOI22V0_8TH40 U849 ( .A1(n41), .A2(n926), .B1(n42), .B2(gpr1_data[23]), .ZN(
        n180) );
  CLKNV1_8TH40 U850 ( .I(n182), .ZN(n926) );
  AOI22V0_8TH40 U851 ( .A1(div_res[54]), .A2(n40), .B1(mul_res_tmp1[54]), .B2(
        n3), .ZN(n185) );
  AOI22V0_8TH40 U852 ( .A1(n41), .A2(n927), .B1(n42), .B2(gpr1_data[22]), .ZN(
        n184) );
  CLKNV1_8TH40 U853 ( .I(n186), .ZN(n927) );
  AOI22V0_8TH40 U854 ( .A1(div_res[53]), .A2(n40), .B1(mul_res_tmp1[53]), .B2(
        n3), .ZN(n188) );
  AOI22V0_8TH40 U855 ( .A1(n41), .A2(n928), .B1(n42), .B2(gpr1_data[21]), .ZN(
        n187) );
  CLKNV1_8TH40 U856 ( .I(n189), .ZN(n928) );
  AOI22V0_8TH40 U857 ( .A1(n41), .A2(n929), .B1(n42), .B2(gpr1_data[20]), .ZN(
        n191) );
  CLKNV1_8TH40 U858 ( .I(n193), .ZN(n929) );
  AOI22V0_8TH40 U859 ( .A1(n41), .A2(n948), .B1(n42), .B2(gpr1_data[1]), .ZN(
        n194) );
  CLKNV1_8TH40 U860 ( .I(n196), .ZN(n948) );
  AOI22V0_8TH40 U861 ( .A1(n41), .A2(n930), .B1(n42), .B2(gpr1_data[19]), .ZN(
        n198) );
  CLKNV1_8TH40 U862 ( .I(n200), .ZN(n930) );
  AOI22V0_8TH40 U863 ( .A1(n41), .A2(n931), .B1(n42), .B2(gpr1_data[18]), .ZN(
        n201) );
  CLKNV1_8TH40 U864 ( .I(n203), .ZN(n931) );
  AOI22V0_8TH40 U865 ( .A1(n41), .A2(n932), .B1(n42), .B2(gpr1_data[17]), .ZN(
        n204) );
  CLKNV1_8TH40 U866 ( .I(n206), .ZN(n932) );
  AOI22V0_8TH40 U867 ( .A1(n41), .A2(n933), .B1(n42), .B2(gpr1_data[16]), .ZN(
        n207) );
  CLKNV1_8TH40 U868 ( .I(n209), .ZN(n933) );
  AOI22V0_8TH40 U869 ( .A1(n41), .A2(n934), .B1(n42), .B2(gpr1_data[15]), .ZN(
        n211) );
  CLKNV1_8TH40 U870 ( .I(n213), .ZN(n934) );
  AOI22V0_8TH40 U871 ( .A1(n41), .A2(n935), .B1(n42), .B2(gpr1_data[14]), .ZN(
        n215) );
  CLKNV1_8TH40 U872 ( .I(n217), .ZN(n935) );
  AOI22V0_8TH40 U873 ( .A1(n41), .A2(n936), .B1(n42), .B2(gpr1_data[13]), .ZN(
        n218) );
  CLKNV1_8TH40 U874 ( .I(n220), .ZN(n936) );
  AOI22V0_8TH40 U875 ( .A1(n41), .A2(n937), .B1(n42), .B2(gpr1_data[12]), .ZN(
        n222) );
  CLKNV1_8TH40 U876 ( .I(n224), .ZN(n937) );
  AOI22V0_8TH40 U877 ( .A1(n41), .A2(n938), .B1(n42), .B2(gpr1_data[11]), .ZN(
        n225) );
  CLKNV1_8TH40 U878 ( .I(n227), .ZN(n938) );
  AOI22V0_8TH40 U879 ( .A1(n41), .A2(n939), .B1(n42), .B2(gpr1_data[10]), .ZN(
        n228) );
  CLKNV1_8TH40 U880 ( .I(n230), .ZN(n939) );
  CLKNV1_8TH40 U881 ( .I(n18), .ZN(n40) );
  AOI22V0_8TH40 U882 ( .A1(n41), .A2(n949), .B1(n42), .B2(gpr1_data[0]), .ZN(
        n232) );
  CLKNV1_8TH40 U883 ( .I(n120), .ZN(n42) );
  NAND3V0P5_8TH40 U884 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n120) );
  CLKNV1_8TH40 U885 ( .I(n237), .ZN(n949) );
  INOR2V0_8TH40 U886 ( .A1(gpr_we), .B1(except_type_o[11]), .ZN(gpr_we_o) );
  OAI21V0_8TH40 U887 ( .A1(n247), .A2(n248), .B(n249), .ZN(n246) );
  AOI222V0_8TH40 U888 ( .A1(mem_cp0_wdata[9]), .A2(n250), .B1(n251), .B2(n972), 
        .C1(N1848), .C2(n252), .ZN(n242) );
  CLKNV1_8TH40 U889 ( .I(n253), .ZN(n972) );
  OAI22V0_8TH40 U890 ( .A1(n28), .A2(n257), .B1(n105), .B2(n258), .ZN(n256) );
  AOI222V0_8TH40 U891 ( .A1(df_memex_lo[9]), .A2(n259), .B1(df_wbex_lo[9]), 
        .B2(n260), .C1(lo_i[9]), .C2(n261), .ZN(n105) );
  AOI222V0_8TH40 U892 ( .A1(df_memex_hi[9]), .A2(n259), .B1(df_wbex_hi[9]), 
        .B2(n260), .C1(hi_i[9]), .C2(n261), .ZN(n28) );
  MUX2NV0_8TH40 U893 ( .I0(n266), .I1(n270), .S(gpr1_data[9]), .ZN(n268) );
  OAI21V0_8TH40 U894 ( .A1(n247), .A2(n276), .B(n249), .ZN(n275) );
  AOI222V0_8TH40 U895 ( .A1(mem_cp0_wdata[8]), .A2(n250), .B1(n251), .B2(n973), 
        .C1(N1847), .C2(n252), .ZN(n273) );
  CLKNV1_8TH40 U896 ( .I(n277), .ZN(n973) );
  OAI22V0_8TH40 U897 ( .A1(n29), .A2(n257), .B1(n106), .B2(n258), .ZN(n278) );
  AOI222V0_8TH40 U898 ( .A1(df_memex_lo[8]), .A2(n259), .B1(df_wbex_lo[8]), 
        .B2(n260), .C1(lo_i[8]), .C2(n261), .ZN(n106) );
  AOI222V0_8TH40 U899 ( .A1(df_memex_hi[8]), .A2(n259), .B1(df_wbex_hi[8]), 
        .B2(n260), .C1(hi_i[8]), .C2(n261), .ZN(n29) );
  MUX2NV0_8TH40 U900 ( .I0(n266), .I1(n270), .S(gpr1_data[8]), .ZN(n281) );
  IOA21V0_8TH40 U901 ( .A1(sum_res[7]), .A2(n244), .B(n249), .ZN(n286) );
  CLKNV1_8TH40 U902 ( .I(n287), .ZN(n974) );
  AO222V0_8TH40 U903 ( .A1(df_memex_lo[7]), .A2(n259), .B1(df_wbex_lo[7]), 
        .B2(n260), .C1(lo_i[7]), .C2(n261), .Z(lo[7]) );
  CLKNV1_8TH40 U904 ( .I(n128), .ZN(n1005) );
  AOI222V0_8TH40 U905 ( .A1(df_memex_hi[7]), .A2(n259), .B1(df_wbex_hi[7]), 
        .B2(n260), .C1(hi_i[7]), .C2(n261), .ZN(n128) );
  MUX2NV0_8TH40 U906 ( .I0(n266), .I1(n270), .S(gpr1_data[7]), .ZN(n292) );
  OAI21V0_8TH40 U907 ( .A1(n298), .A2(n299), .B(n300), .ZN(n297) );
  CLKNV1_8TH40 U908 ( .I(n301), .ZN(n975) );
  OAI22V0_8TH40 U909 ( .A1(n30), .A2(n257), .B1(n107), .B2(n258), .ZN(n302) );
  AOI222V0_8TH40 U910 ( .A1(df_memex_lo[6]), .A2(n259), .B1(df_wbex_lo[6]), 
        .B2(n260), .C1(lo_i[6]), .C2(n261), .ZN(n107) );
  AOI222V0_8TH40 U911 ( .A1(df_memex_hi[6]), .A2(n259), .B1(df_wbex_hi[6]), 
        .B2(n260), .C1(hi_i[6]), .C2(n261), .ZN(n30) );
  MUX2NV0_8TH40 U912 ( .I0(n266), .I1(n270), .S(gpr1_data[6]), .ZN(n305) );
  MUX2NV0_8TH40 U913 ( .I0(n317), .I1(n321), .S(gpr1_data[5]), .ZN(n320) );
  MUX2NV0_8TH40 U914 ( .I0(n322), .I1(n323), .S(gpr1_data[1]), .ZN(n312) );
  NAND3V0P5_8TH40 U915 ( .A1(n324), .A2(gpr1_data[0]), .A3(n325), .ZN(n323) );
  NAND3V0P5_8TH40 U916 ( .A1(n326), .A2(n912), .A3(n327), .ZN(n322) );
  CLKNV1_8TH40 U917 ( .I(n135), .ZN(n1007) );
  AOI222V0_8TH40 U918 ( .A1(df_memex_hi[5]), .A2(n259), .B1(df_wbex_hi[5]), 
        .B2(n260), .C1(hi_i[5]), .C2(n261), .ZN(n135) );
  AO222V0_8TH40 U919 ( .A1(df_memex_lo[5]), .A2(n259), .B1(df_wbex_lo[5]), 
        .B2(n260), .C1(lo_i[5]), .C2(n261), .Z(lo[5]) );
  AOI22V0_8TH40 U920 ( .A1(link_addr[5]), .A2(n245), .B1(n251), .B2(n976), 
        .ZN(n306) );
  CLKNV1_8TH40 U921 ( .I(n330), .ZN(n976) );
  MUX2NV0_8TH40 U922 ( .I0(n266), .I1(n270), .S(gpr1_data[4]), .ZN(n340) );
  AOI222V0_8TH40 U923 ( .A1(df_memex_hi[4]), .A2(n259), .B1(df_wbex_hi[4]), 
        .B2(n260), .C1(hi_i[4]), .C2(n261), .ZN(n31) );
  AOI222V0_8TH40 U924 ( .A1(df_memex_lo[4]), .A2(n259), .B1(df_wbex_lo[4]), 
        .B2(n260), .C1(lo_i[4]), .C2(n261), .ZN(n108) );
  CLKNAND2V1_8TH40 U925 ( .A1(gpr1_data[7]), .A2(gpr1_data[9]), .ZN(n349) );
  CLKNV1_8TH40 U926 ( .I(n350), .ZN(n347) );
  OAOI211V0_8TH40 U927 ( .A1(n1033), .A2(n1035), .B(n351), .C(n352), .ZN(n344)
         );
  INAND3V0_8TH40 U928 ( .A1(n359), .B1(n1030), .B2(gpr1_data[15]), .ZN(n357)
         );
  OAOI211V0_8TH40 U929 ( .A1(gpr1_data[13]), .A2(gpr1_data[11]), .B(n360), .C(
        n361), .ZN(n355) );
  AOI22V0_8TH40 U930 ( .A1(link_addr[4]), .A2(n245), .B1(n251), .B2(n977), 
        .ZN(n332) );
  CLKNV1_8TH40 U931 ( .I(n362), .ZN(n977) );
  OAI22V0_8TH40 U932 ( .A1(n1029), .A2(n376), .B1(n377), .B2(n378), .ZN(n375)
         );
  OAI221V0_8TH40 U933 ( .A1(n1023), .A2(n379), .B1(n1040), .B2(n380), .C(n381), 
        .ZN(n373) );
  CLKNV1_8TH40 U934 ( .I(n382), .ZN(n380) );
  AOAI211V0_8TH40 U935 ( .A1(gpr1_data[19]), .A2(gpr1_data[21]), .B(n386), .C(
        n387), .ZN(n385) );
  OAI211V0_8TH40 U936 ( .A1(gpr1_data[7]), .A2(n388), .B(n389), .C(n390), .ZN(
        n384) );
  CLKNV1_8TH40 U937 ( .I(n391), .ZN(n978) );
  AOI22V0_8TH40 U938 ( .A1(mem_cp0_wdata[3]), .A2(n250), .B1(n288), .B2(lo[3]), 
        .ZN(n367) );
  AO222V0_8TH40 U939 ( .A1(df_memex_lo[3]), .A2(n259), .B1(df_wbex_lo[3]), 
        .B2(n260), .C1(lo_i[3]), .C2(n261), .Z(lo[3]) );
  OR2V0_8TH40 U940 ( .A1(n249), .A2(N1873), .Z(n300) );
  AOI221V0_8TH40 U941 ( .A1(n325), .A2(n913), .B1(n395), .B2(n396), .C(n397), 
        .ZN(n394) );
  CLKNV1_8TH40 U942 ( .I(n400), .ZN(n399) );
  OAI22V0_8TH40 U943 ( .A1(n913), .A2(n401), .B1(n402), .B2(n403), .ZN(n398)
         );
  MUX2NV0_8TH40 U944 ( .I0(n266), .I1(n270), .S(gpr1_data[3]), .ZN(n405) );
  CLKNV1_8TH40 U945 ( .I(n142), .ZN(n1009) );
  AOI222V0_8TH40 U946 ( .A1(df_memex_hi[3]), .A2(n259), .B1(df_wbex_hi[3]), 
        .B2(n260), .C1(hi_i[3]), .C2(n261), .ZN(n142) );
  MUX2NV0_8TH40 U947 ( .I0(n413), .I1(n314), .S(gpr1_data[31]), .ZN(n412) );
  CLKNAND2V1_8TH40 U948 ( .A1(n265), .A2(n1042), .ZN(n413) );
  AO211V0_8TH40 U949 ( .A1(gpr1_data[31]), .A2(n270), .B(n319), .C(n416), .Z(
        n415) );
  AOI222V0_8TH40 U950 ( .A1(n289), .A2(n981), .B1(mem_cp0_wdata[31]), .B2(n250), .C1(n288), .C2(lo[31]), .ZN(n408) );
  AO222V0_8TH40 U951 ( .A1(df_memex_lo[31]), .A2(n259), .B1(df_wbex_lo[31]), 
        .B2(n260), .C1(lo_i[31]), .C2(n261), .Z(lo[31]) );
  CLKNV1_8TH40 U952 ( .I(n146), .ZN(n981) );
  AOI222V0_8TH40 U953 ( .A1(df_memex_hi[31]), .A2(n259), .B1(df_wbex_hi[31]), 
        .B2(n260), .C1(hi_i[31]), .C2(n261), .ZN(n146) );
  AOI22V0_8TH40 U954 ( .A1(n244), .A2(sum_res[31]), .B1(link_addr[31]), .B2(
        n245), .ZN(n407) );
  CLKNV1_8TH40 U955 ( .I(n417), .ZN(n950) );
  IOA21V0_8TH40 U956 ( .A1(n423), .A2(n416), .B(n424), .ZN(n422) );
  CLKNV1_8TH40 U957 ( .I(n425), .ZN(n951) );
  OAI22V0_8TH40 U958 ( .A1(n19), .A2(n257), .B1(n109), .B2(n258), .ZN(n426) );
  AOI222V0_8TH40 U959 ( .A1(df_memex_lo[30]), .A2(n259), .B1(df_wbex_lo[30]), 
        .B2(n260), .C1(lo_i[30]), .C2(n261), .ZN(n109) );
  AOI222V0_8TH40 U960 ( .A1(df_memex_hi[30]), .A2(n259), .B1(df_wbex_hi[30]), 
        .B2(n260), .C1(hi_i[30]), .C2(n261), .ZN(n19) );
  MUX2NV0_8TH40 U961 ( .I0(n266), .I1(n270), .S(gpr1_data[30]), .ZN(n429) );
  OAI22V0_8TH40 U962 ( .A1(n32), .A2(n257), .B1(n110), .B2(n258), .ZN(n434) );
  AOI222V0_8TH40 U963 ( .A1(df_memex_lo[2]), .A2(n259), .B1(df_wbex_lo[2]), 
        .B2(n260), .C1(lo_i[2]), .C2(n261), .ZN(n110) );
  AOI222V0_8TH40 U964 ( .A1(df_memex_hi[2]), .A2(n259), .B1(df_wbex_hi[2]), 
        .B2(n260), .C1(hi_i[2]), .C2(n261), .ZN(n32) );
  MUX2NV0_8TH40 U965 ( .I0(n317), .I1(n321), .S(gpr1_data[2]), .ZN(n436) );
  AOI221V0_8TH40 U966 ( .A1(n446), .A2(n447), .B1(n448), .B2(gpr1_data[18]), 
        .C(n449), .ZN(n445) );
  CLKNV1_8TH40 U967 ( .I(n454), .ZN(n453) );
  NAND4V0P5_8TH40 U968 ( .A1(n455), .A2(gpr1_data[3]), .A3(n916), .A4(n1041), 
        .ZN(n443) );
  AOI221V0_8TH40 U969 ( .A1(n461), .A2(n462), .B1(n348), .B2(n1036), .C(n463), 
        .ZN(n460) );
  AOI21V0_8TH40 U970 ( .A1(gpr1_data[26]), .A2(gpr1_data[27]), .B(n467), .ZN(
        n466) );
  NAND4V0P5_8TH40 U971 ( .A1(n395), .A2(gpr1_data[5]), .A3(gpr1_data[4]), .A4(
        n915), .ZN(n457) );
  AOI22V0_8TH40 U972 ( .A1(link_addr[2]), .A2(n245), .B1(n251), .B2(n979), 
        .ZN(n438) );
  CLKNV1_8TH40 U973 ( .I(n468), .ZN(n979) );
  MUX2NV0_8TH40 U974 ( .I0(n317), .I1(n321), .S(gpr1_data[29]), .ZN(n479) );
  CLKNV1_8TH40 U975 ( .I(n156), .ZN(n983) );
  AOI222V0_8TH40 U976 ( .A1(df_memex_hi[29]), .A2(n259), .B1(df_wbex_hi[29]), 
        .B2(n260), .C1(hi_i[29]), .C2(n261), .ZN(n156) );
  AO222V0_8TH40 U977 ( .A1(df_memex_lo[29]), .A2(n259), .B1(df_wbex_lo[29]), 
        .B2(n260), .C1(lo_i[29]), .C2(n261), .Z(lo[29]) );
  CLKNV1_8TH40 U978 ( .I(n480), .ZN(n329) );
  AOI22V0_8TH40 U979 ( .A1(link_addr[29]), .A2(n245), .B1(n251), .B2(n952), 
        .ZN(n469) );
  CLKNV1_8TH40 U980 ( .I(n481), .ZN(n952) );
  IOA21V0_8TH40 U981 ( .A1(n487), .A2(n416), .B(n424), .ZN(n486) );
  CLKNV1_8TH40 U982 ( .I(n488), .ZN(n953) );
  OAI22V0_8TH40 U983 ( .A1(n20), .A2(n257), .B1(n111), .B2(n258), .ZN(n489) );
  AOI222V0_8TH40 U984 ( .A1(df_memex_lo[28]), .A2(n259), .B1(df_wbex_lo[28]), 
        .B2(n260), .C1(lo_i[28]), .C2(n261), .ZN(n111) );
  AOI222V0_8TH40 U985 ( .A1(df_memex_hi[28]), .A2(n259), .B1(df_wbex_hi[28]), 
        .B2(n260), .C1(hi_i[28]), .C2(n261), .ZN(n20) );
  MUX2NV0_8TH40 U986 ( .I0(n266), .I1(n270), .S(gpr1_data[28]), .ZN(n492) );
  MUX2NV0_8TH40 U987 ( .I0(n317), .I1(n321), .S(gpr1_data[27]), .ZN(n502) );
  CLKNV1_8TH40 U988 ( .I(n163), .ZN(n985) );
  AOI222V0_8TH40 U989 ( .A1(df_memex_hi[27]), .A2(n259), .B1(df_wbex_hi[27]), 
        .B2(n260), .C1(hi_i[27]), .C2(n261), .ZN(n163) );
  AO222V0_8TH40 U990 ( .A1(df_memex_lo[27]), .A2(n259), .B1(df_wbex_lo[27]), 
        .B2(n260), .C1(lo_i[27]), .C2(n261), .Z(lo[27]) );
  AOI22V0_8TH40 U991 ( .A1(link_addr[27]), .A2(n245), .B1(n251), .B2(n954), 
        .ZN(n493) );
  CLKNV1_8TH40 U992 ( .I(n504), .ZN(n954) );
  MUX2NV0_8TH40 U993 ( .I0(n317), .I1(n321), .S(gpr1_data[26]), .ZN(n514) );
  CLKNV1_8TH40 U994 ( .I(n167), .ZN(n986) );
  AOI222V0_8TH40 U995 ( .A1(df_memex_hi[26]), .A2(n259), .B1(df_wbex_hi[26]), 
        .B2(n260), .C1(hi_i[26]), .C2(n261), .ZN(n167) );
  AO222V0_8TH40 U996 ( .A1(df_memex_lo[26]), .A2(n259), .B1(df_wbex_lo[26]), 
        .B2(n260), .C1(lo_i[26]), .C2(n261), .Z(lo[26]) );
  AOI22V0_8TH40 U997 ( .A1(link_addr[26]), .A2(n245), .B1(n251), .B2(n955), 
        .ZN(n505) );
  CLKNV1_8TH40 U998 ( .I(n515), .ZN(n955) );
  MUX2NV0_8TH40 U999 ( .I0(n317), .I1(n321), .S(gpr1_data[25]), .ZN(n525) );
  CLKNV1_8TH40 U1000 ( .I(n171), .ZN(n987) );
  AOI222V0_8TH40 U1001 ( .A1(df_memex_hi[25]), .A2(n259), .B1(df_wbex_hi[25]), 
        .B2(n260), .C1(hi_i[25]), .C2(n261), .ZN(n171) );
  AO222V0_8TH40 U1002 ( .A1(df_memex_lo[25]), .A2(n259), .B1(df_wbex_lo[25]), 
        .B2(n260), .C1(lo_i[25]), .C2(n261), .Z(lo[25]) );
  AOI22V0_8TH40 U1003 ( .A1(link_addr[25]), .A2(n245), .B1(n251), .B2(n956), 
        .ZN(n516) );
  CLKNV1_8TH40 U1004 ( .I(n527), .ZN(n956) );
  MUX2NV0_8TH40 U1005 ( .I0(n317), .I1(n321), .S(gpr1_data[24]), .ZN(n537) );
  CLKNV1_8TH40 U1006 ( .I(n538), .ZN(n476) );
  CLKNV1_8TH40 U1007 ( .I(n175), .ZN(n988) );
  AOI222V0_8TH40 U1008 ( .A1(df_memex_hi[24]), .A2(n259), .B1(df_wbex_hi[24]), 
        .B2(n260), .C1(hi_i[24]), .C2(n261), .ZN(n175) );
  AO222V0_8TH40 U1009 ( .A1(df_memex_lo[24]), .A2(n259), .B1(df_wbex_lo[24]), 
        .B2(n260), .C1(lo_i[24]), .C2(n261), .Z(lo[24]) );
  AOI22V0_8TH40 U1010 ( .A1(link_addr[24]), .A2(n245), .B1(n251), .B2(n957), 
        .ZN(n528) );
  CLKNV1_8TH40 U1011 ( .I(n540), .ZN(n957) );
  CLKNV1_8TH40 U1012 ( .I(n546), .ZN(n958) );
  AOI222V0_8TH40 U1013 ( .A1(n289), .A2(n989), .B1(mem_cp0_wdata[23]), .B2(
        n250), .C1(n288), .C2(lo[23]), .ZN(n543) );
  AO222V0_8TH40 U1014 ( .A1(df_memex_lo[23]), .A2(n259), .B1(df_wbex_lo[23]), 
        .B2(n260), .C1(lo_i[23]), .C2(n261), .Z(lo[23]) );
  CLKNV1_8TH40 U1015 ( .I(n179), .ZN(n989) );
  AOI222V0_8TH40 U1016 ( .A1(df_memex_hi[23]), .A2(n259), .B1(df_wbex_hi[23]), 
        .B2(n260), .C1(hi_i[23]), .C2(n261), .ZN(n179) );
  OAI21V0_8TH40 U1017 ( .A1(n1042), .A2(n548), .B(n424), .ZN(n538) );
  MUX2NV0_8TH40 U1018 ( .I0(n266), .I1(n270), .S(gpr1_data[23]), .ZN(n550) );
  MUX2NV0_8TH40 U1019 ( .I0(n317), .I1(n321), .S(gpr1_data[22]), .ZN(n561) );
  CLKNV1_8TH40 U1020 ( .I(n183), .ZN(n990) );
  AOI222V0_8TH40 U1021 ( .A1(df_memex_hi[22]), .A2(n259), .B1(df_wbex_hi[22]), 
        .B2(n260), .C1(hi_i[22]), .C2(n261), .ZN(n183) );
  AO222V0_8TH40 U1022 ( .A1(df_memex_lo[22]), .A2(n259), .B1(df_wbex_lo[22]), 
        .B2(n260), .C1(lo_i[22]), .C2(n261), .Z(lo[22]) );
  AOI22V0_8TH40 U1023 ( .A1(link_addr[22]), .A2(n245), .B1(n251), .B2(n959), 
        .ZN(n551) );
  CLKNV1_8TH40 U1024 ( .I(n562), .ZN(n959) );
  OAI21V0_8TH40 U1025 ( .A1(n480), .A2(n548), .B(n424), .ZN(n567) );
  CLKNV1_8TH40 U1026 ( .I(n568), .ZN(n960) );
  OAI22V0_8TH40 U1027 ( .A1(n21), .A2(n257), .B1(n112), .B2(n258), .ZN(n569)
         );
  AOI222V0_8TH40 U1028 ( .A1(df_memex_lo[21]), .A2(n259), .B1(df_wbex_lo[21]), 
        .B2(n260), .C1(lo_i[21]), .C2(n261), .ZN(n112) );
  AOI222V0_8TH40 U1029 ( .A1(df_memex_hi[21]), .A2(n259), .B1(df_wbex_hi[21]), 
        .B2(n260), .C1(hi_i[21]), .C2(n261), .ZN(n21) );
  MUX2NV0_8TH40 U1030 ( .I0(n266), .I1(n270), .S(gpr1_data[21]), .ZN(n572) );
  MUX2NV0_8TH40 U1031 ( .I0(n317), .I1(n321), .S(gpr1_data[20]), .ZN(n582) );
  CLKNV1_8TH40 U1032 ( .I(n583), .ZN(n558) );
  CLKNV1_8TH40 U1033 ( .I(n190), .ZN(n992) );
  AOI222V0_8TH40 U1034 ( .A1(df_memex_hi[20]), .A2(n259), .B1(df_wbex_hi[20]), 
        .B2(n260), .C1(hi_i[20]), .C2(n261), .ZN(n190) );
  AO222V0_8TH40 U1035 ( .A1(df_memex_lo[20]), .A2(n259), .B1(df_wbex_lo[20]), 
        .B2(n260), .C1(lo_i[20]), .C2(n261), .Z(lo[20]) );
  AOI22V0_8TH40 U1036 ( .A1(link_addr[20]), .A2(n245), .B1(n251), .B2(n961), 
        .ZN(n573) );
  CLKNV1_8TH40 U1037 ( .I(n584), .ZN(n961) );
  OAI22V0_8TH40 U1038 ( .A1(n33), .A2(n257), .B1(n113), .B2(n258), .ZN(n589)
         );
  AOI222V0_8TH40 U1039 ( .A1(df_memex_lo[1]), .A2(n259), .B1(df_wbex_lo[1]), 
        .B2(n260), .C1(lo_i[1]), .C2(n261), .ZN(n113) );
  AOI222V0_8TH40 U1040 ( .A1(df_memex_hi[1]), .A2(n259), .B1(df_wbex_hi[1]), 
        .B2(n260), .C1(hi_i[1]), .C2(n261), .ZN(n33) );
  MUX2NV0_8TH40 U1041 ( .I0(n317), .I1(n321), .S(gpr1_data[1]), .ZN(n591) );
  OAI31V0_8TH40 U1042 ( .A1(n376), .A2(gpr1_data[18]), .A3(n1029), .B(n356), 
        .ZN(n605) );
  NAND3V0P5_8TH40 U1043 ( .A1(n606), .A2(gpr1_data[9]), .A3(n446), .ZN(n356)
         );
  NOR2V0P5_8TH40 U1044 ( .A1(n1038), .A2(n609), .ZN(n608) );
  OAI22V0_8TH40 U1045 ( .A1(n1041), .A2(n403), .B1(n451), .B2(n454), .ZN(n602)
         );
  CLKNV1_8TH40 U1046 ( .I(n610), .ZN(n601) );
  AOI33V0_8TH40 U1047 ( .A1(gpr1_data[13]), .A2(n1032), .A3(n360), .B1(
        gpr1_data[21]), .B2(n1024), .B3(n611), .ZN(n599) );
  CLKNV1_8TH40 U1048 ( .I(n299), .ZN(n328) );
  AOI31V0_8TH40 U1049 ( .A1(gpr1_data[30]), .A2(gpr1_data[31]), .A3(n616), .B(
        n617), .ZN(n615) );
  AOI22V0_8TH40 U1050 ( .A1(n395), .A2(n1041), .B1(n618), .B2(n1026), .ZN(n614) );
  OAI31V0_8TH40 U1051 ( .A1(n622), .A2(n1036), .A3(n623), .B(n387), .ZN(n621)
         );
  NAND3V0P5_8TH40 U1052 ( .A1(n624), .A2(n1029), .A3(n461), .ZN(n387) );
  OAI21V0_8TH40 U1053 ( .A1(n1021), .A2(n1022), .B(n625), .ZN(n619) );
  OAI32V0_8TH40 U1054 ( .A1(n1024), .A2(gpr1_data[21]), .A3(n386), .B1(n626), 
        .B2(n464), .ZN(n613) );
  CLKNV1_8TH40 U1055 ( .I(n346), .ZN(n324) );
  AOI22V0_8TH40 U1056 ( .A1(link_addr[1]), .A2(n245), .B1(n251), .B2(n980), 
        .ZN(n593) );
  CLKNV1_8TH40 U1057 ( .I(n627), .ZN(n980) );
  CLKNV1_8TH40 U1058 ( .I(n633), .ZN(n962) );
  AOI222V0_8TH40 U1059 ( .A1(n289), .A2(n993), .B1(mem_cp0_wdata[19]), .B2(
        n250), .C1(n288), .C2(lo[19]), .ZN(n630) );
  AO222V0_8TH40 U1060 ( .A1(df_memex_lo[19]), .A2(n259), .B1(df_wbex_lo[19]), 
        .B2(n260), .C1(lo_i[19]), .C2(n261), .Z(lo[19]) );
  CLKNV1_8TH40 U1061 ( .I(n197), .ZN(n993) );
  AOI222V0_8TH40 U1062 ( .A1(df_memex_hi[19]), .A2(n259), .B1(df_wbex_hi[19]), 
        .B2(n260), .C1(hi_i[19]), .C2(n261), .ZN(n197) );
  OAI21V0_8TH40 U1063 ( .A1(n635), .A2(n548), .B(n424), .ZN(n583) );
  CLKNV1_8TH40 U1064 ( .I(n503), .ZN(n635) );
  MUX2NV0_8TH40 U1065 ( .I0(n266), .I1(n270), .S(gpr1_data[19]), .ZN(n637) );
  OAI21V0_8TH40 U1066 ( .A1(n643), .A2(n548), .B(n424), .ZN(n642) );
  CLKNV1_8TH40 U1067 ( .I(n644), .ZN(n963) );
  OAI22V0_8TH40 U1068 ( .A1(n22), .A2(n257), .B1(n114), .B2(n258), .ZN(n645)
         );
  AOI222V0_8TH40 U1069 ( .A1(df_memex_lo[18]), .A2(n259), .B1(df_wbex_lo[18]), 
        .B2(n260), .C1(lo_i[18]), .C2(n261), .ZN(n114) );
  AOI222V0_8TH40 U1070 ( .A1(df_memex_hi[18]), .A2(n259), .B1(df_wbex_hi[18]), 
        .B2(n260), .C1(hi_i[18]), .C2(n261), .ZN(n22) );
  MUX2NV0_8TH40 U1071 ( .I0(n266), .I1(n270), .S(gpr1_data[18]), .ZN(n648) );
  OAI21V0_8TH40 U1072 ( .A1(n248), .A2(n548), .B(n424), .ZN(n653) );
  CLKNV1_8TH40 U1073 ( .I(n526), .ZN(n248) );
  INOR2V0_8TH40 U1074 ( .A1(n503), .B1(N1872), .ZN(n526) );
  CLKNV1_8TH40 U1075 ( .I(n654), .ZN(n964) );
  OAI22V0_8TH40 U1076 ( .A1(n23), .A2(n257), .B1(n115), .B2(n258), .ZN(n655)
         );
  AOI222V0_8TH40 U1077 ( .A1(df_memex_lo[17]), .A2(n259), .B1(df_wbex_lo[17]), 
        .B2(n260), .C1(lo_i[17]), .C2(n261), .ZN(n115) );
  AOI222V0_8TH40 U1078 ( .A1(df_memex_hi[17]), .A2(n259), .B1(df_wbex_hi[17]), 
        .B2(n260), .C1(hi_i[17]), .C2(n261), .ZN(n23) );
  MUX2NV0_8TH40 U1079 ( .I0(n266), .I1(n270), .S(gpr1_data[17]), .ZN(n658) );
  OAI21V0_8TH40 U1080 ( .A1(n276), .A2(n548), .B(n424), .ZN(n663) );
  CLKNAND2V1_8TH40 U1081 ( .A1(n416), .A2(n2), .ZN(n548) );
  NOR2V0P5_8TH40 U1082 ( .A1(n664), .A2(n17), .ZN(n416) );
  CLKNV1_8TH40 U1083 ( .I(n665), .ZN(n965) );
  OAI22V0_8TH40 U1084 ( .A1(n24), .A2(n257), .B1(n116), .B2(n258), .ZN(n666)
         );
  AOI222V0_8TH40 U1085 ( .A1(df_memex_lo[16]), .A2(n259), .B1(df_wbex_lo[16]), 
        .B2(n260), .C1(lo_i[16]), .C2(n261), .ZN(n116) );
  AOI222V0_8TH40 U1086 ( .A1(df_memex_hi[16]), .A2(n259), .B1(df_wbex_hi[16]), 
        .B2(n260), .C1(hi_i[16]), .C2(n261), .ZN(n24) );
  MUX2NV0_8TH40 U1087 ( .I0(n266), .I1(n270), .S(gpr1_data[16]), .ZN(n669) );
  IOA21V0_8TH40 U1088 ( .A1(sum_res[15]), .A2(n244), .B(n424), .ZN(n674) );
  CLKNV1_8TH40 U1089 ( .I(n675), .ZN(n966) );
  AO222V0_8TH40 U1090 ( .A1(df_memex_lo[15]), .A2(n259), .B1(df_wbex_lo[15]), 
        .B2(n260), .C1(lo_i[15]), .C2(n261), .Z(lo[15]) );
  CLKNV1_8TH40 U1091 ( .I(n210), .ZN(n997) );
  AOI222V0_8TH40 U1092 ( .A1(df_memex_hi[15]), .A2(n259), .B1(df_wbex_hi[15]), 
        .B2(n260), .C1(hi_i[15]), .C2(n261), .ZN(n210) );
  MUX2NV0_8TH40 U1093 ( .I0(n266), .I1(n270), .S(gpr1_data[15]), .ZN(n678) );
  MUX2NV0_8TH40 U1094 ( .I0(n266), .I1(n270), .S(gpr1_data[14]), .ZN(n687) );
  CLKNV1_8TH40 U1095 ( .I(n214), .ZN(n998) );
  AOI222V0_8TH40 U1096 ( .A1(df_memex_hi[14]), .A2(n259), .B1(df_wbex_hi[14]), 
        .B2(n260), .C1(hi_i[14]), .C2(n261), .ZN(n214) );
  AO222V0_8TH40 U1097 ( .A1(df_memex_lo[14]), .A2(n259), .B1(df_wbex_lo[14]), 
        .B2(n260), .C1(lo_i[14]), .C2(n261), .Z(lo[14]) );
  CLKNAND2V1_8TH40 U1098 ( .A1(n298), .A2(n689), .ZN(n423) );
  AOI22V0_8TH40 U1099 ( .A1(link_addr[14]), .A2(n245), .B1(n251), .B2(n967), 
        .ZN(n679) );
  CLKNV1_8TH40 U1100 ( .I(n690), .ZN(n967) );
  OAI21V0_8TH40 U1101 ( .A1(n480), .A2(n247), .B(n249), .ZN(n695) );
  NOR2V0P5_8TH40 U1102 ( .A1(n503), .A2(n696), .ZN(n480) );
  CLKNV1_8TH40 U1103 ( .I(n697), .ZN(n968) );
  OAI22V0_8TH40 U1104 ( .A1(n25), .A2(n257), .B1(n117), .B2(n258), .ZN(n698)
         );
  AOI222V0_8TH40 U1105 ( .A1(df_memex_lo[13]), .A2(n259), .B1(df_wbex_lo[13]), 
        .B2(n260), .C1(lo_i[13]), .C2(n261), .ZN(n117) );
  AOI222V0_8TH40 U1106 ( .A1(df_memex_hi[13]), .A2(n259), .B1(df_wbex_hi[13]), 
        .B2(n260), .C1(hi_i[13]), .C2(n261), .ZN(n25) );
  MUX2NV0_8TH40 U1107 ( .I0(n266), .I1(n270), .S(gpr1_data[13]), .ZN(n701) );
  MUX2NV0_8TH40 U1108 ( .I0(n266), .I1(n270), .S(gpr1_data[12]), .ZN(n710) );
  CLKNV1_8TH40 U1109 ( .I(n221), .ZN(n1000) );
  AOI222V0_8TH40 U1110 ( .A1(df_memex_hi[12]), .A2(n259), .B1(df_wbex_hi[12]), 
        .B2(n260), .C1(hi_i[12]), .C2(n261), .ZN(n221) );
  AO222V0_8TH40 U1111 ( .A1(df_memex_lo[12]), .A2(n259), .B1(df_wbex_lo[12]), 
        .B2(n260), .C1(lo_i[12]), .C2(n261), .Z(lo[12]) );
  CLKNAND2V1_8TH40 U1112 ( .A1(n689), .A2(n353), .ZN(n487) );
  AOI21V0_8TH40 U1113 ( .A1(n2), .A2(gpr2_data[31]), .B(n503), .ZN(n689) );
  NOR2V0P5_8TH40 U1114 ( .A1(n1042), .A2(N1873), .ZN(n503) );
  AOI22V0_8TH40 U1115 ( .A1(link_addr[12]), .A2(n245), .B1(n251), .B2(n969), 
        .ZN(n702) );
  CLKNV1_8TH40 U1116 ( .I(n711), .ZN(n969) );
  OAI21V0_8TH40 U1117 ( .A1(N1873), .A2(n424), .B(n249), .ZN(n716) );
  AOI222V0_8TH40 U1118 ( .A1(mem_cp0_wdata[11]), .A2(n250), .B1(n251), .B2(
        n970), .C1(N1850), .C2(n252), .ZN(n714) );
  CLKNV1_8TH40 U1119 ( .I(n717), .ZN(n970) );
  OAI22V0_8TH40 U1120 ( .A1(n26), .A2(n257), .B1(n118), .B2(n258), .ZN(n718)
         );
  AOI222V0_8TH40 U1121 ( .A1(df_memex_lo[11]), .A2(n259), .B1(df_wbex_lo[11]), 
        .B2(n260), .C1(lo_i[11]), .C2(n261), .ZN(n118) );
  AOI222V0_8TH40 U1122 ( .A1(df_memex_hi[11]), .A2(n259), .B1(df_wbex_hi[11]), 
        .B2(n260), .C1(hi_i[11]), .C2(n261), .ZN(n26) );
  MUX2NV0_8TH40 U1123 ( .I0(n266), .I1(n270), .S(gpr1_data[11]), .ZN(n721) );
  OAI21V0_8TH40 U1124 ( .A1(n247), .A2(n643), .B(n249), .ZN(n726) );
  CLKNAND2V1_8TH40 U1125 ( .A1(n727), .A2(n2), .ZN(n249) );
  CLKNV1_8TH40 U1126 ( .I(n424), .ZN(n727) );
  CLKNAND2V1_8TH40 U1127 ( .A1(n688), .A2(gpr2_data[31]), .ZN(n424) );
  CLKNV1_8TH40 U1128 ( .I(n441), .ZN(n643) );
  NOR2V0P5_8TH40 U1129 ( .A1(n298), .A2(N1873), .ZN(n441) );
  AOI21V0_8TH40 U1130 ( .A1(n912), .A2(gpr2_data[31]), .B(n696), .ZN(n298) );
  CLKNV1_8TH40 U1131 ( .I(n688), .ZN(n247) );
  AOI222V0_8TH40 U1132 ( .A1(mem_cp0_wdata[10]), .A2(n250), .B1(n251), .B2(
        n971), .C1(N1849), .C2(n252), .ZN(n724) );
  CLKNV1_8TH40 U1133 ( .I(n728), .ZN(n971) );
  OAI22V0_8TH40 U1134 ( .A1(n27), .A2(n257), .B1(n119), .B2(n258), .ZN(n729)
         );
  AOI222V0_8TH40 U1135 ( .A1(df_memex_lo[10]), .A2(n259), .B1(df_wbex_lo[10]), 
        .B2(n260), .C1(lo_i[10]), .C2(n261), .ZN(n119) );
  AOI222V0_8TH40 U1136 ( .A1(df_memex_hi[10]), .A2(n259), .B1(df_wbex_hi[10]), 
        .B2(n260), .C1(hi_i[10]), .C2(n261), .ZN(n27) );
  MUX2NV0_8TH40 U1137 ( .I0(n266), .I1(n270), .S(gpr1_data[10]), .ZN(n732) );
  CLKNV1_8TH40 U1138 ( .I(n321), .ZN(n270) );
  CLKNV1_8TH40 U1139 ( .I(n317), .ZN(n266) );
  CLKNV1_8TH40 U1140 ( .I(n316), .ZN(n265) );
  NOR4V0P5_8TH40 U1141 ( .A1(n745), .A2(n746), .A3(n747), .A4(n748), .ZN(n744)
         );
  I2NOR3V1_8TH40 U1142 ( .A1(n749), .A2(n750), .B(n751), .ZN(n255) );
  MUX2NV0_8TH40 U1143 ( .I0(n317), .I1(n321), .S(gpr1_data[0]), .ZN(n753) );
  CLKNAND2V1_8TH40 U1144 ( .A1(n754), .A2(n742), .ZN(n321) );
  CLKNV1_8TH40 U1145 ( .I(n269), .ZN(n319) );
  CLKNAND2V1_8TH40 U1146 ( .A1(n754), .A2(n755), .ZN(n317) );
  NAND3V0P5_8TH40 U1147 ( .A1(inst_type[0]), .A2(inst_type[1]), .A3(n754), 
        .ZN(n316) );
  CLKNV1_8TH40 U1148 ( .I(n263), .ZN(n314) );
  NAND4V0P5_8TH40 U1149 ( .A1(n757), .A2(n758), .A3(n759), .A4(n235), .ZN(n756) );
  CLKNAND2V1_8TH40 U1150 ( .A1(n754), .A2(n236), .ZN(n269) );
  NOR3V0P5_8TH40 U1151 ( .A1(inst_class[1]), .A2(rst), .A3(inst_class[2]), 
        .ZN(n761) );
  AOI22V0_8TH40 U1152 ( .A1(mem_cp0_wdata[0]), .A2(n250), .B1(n288), .B2(lo[0]), .ZN(n738) );
  AO222V0_8TH40 U1153 ( .A1(df_memex_lo[0]), .A2(n259), .B1(df_wbex_lo[0]), 
        .B2(n260), .C1(lo_i[0]), .C2(n261), .Z(lo[0]) );
  CLKNV1_8TH40 U1154 ( .I(n258), .ZN(n288) );
  NAND4V0P5_8TH40 U1155 ( .A1(n757), .A2(n755), .A3(n234), .A4(n764), .ZN(n258) );
  INOR2V0_8TH40 U1156 ( .A1(n749), .B1(n750), .ZN(n250) );
  AND3V0_8TH40 U1157 ( .A1(n751), .A2(n750), .A3(n749), .Z(n254) );
  AND2V0_8TH40 U1158 ( .A1(N2186), .A2(n757), .Z(n749) );
  CLKXOR2V2_8TH40 U1159 ( .A1(mem_cp0_waddr[2]), .A2(inst_i[13]), .Z(n770) );
  CLKXOR2V2_8TH40 U1160 ( .A1(mem_cp0_waddr[4]), .A2(inst_i[15]), .Z(n769) );
  CLKXOR2V2_8TH40 U1161 ( .A1(mem_cp0_waddr[3]), .A2(inst_i[14]), .Z(n768) );
  XNOR2V0_8TH40 U1162 ( .A1(inst_i[11]), .A2(mem_cp0_waddr[0]), .ZN(n766) );
  XNOR2V0_8TH40 U1163 ( .A1(inst_i[12]), .A2(mem_cp0_waddr[1]), .ZN(n765) );
  CLKXOR2V2_8TH40 U1164 ( .A1(wb_cp0_waddr[2]), .A2(inst_i[13]), .Z(n776) );
  CLKXOR2V2_8TH40 U1165 ( .A1(wb_cp0_waddr[4]), .A2(inst_i[15]), .Z(n775) );
  CLKXOR2V2_8TH40 U1166 ( .A1(wb_cp0_waddr[3]), .A2(inst_i[14]), .Z(n774) );
  XNOR2V0_8TH40 U1167 ( .A1(inst_i[11]), .A2(wb_cp0_waddr[0]), .ZN(n772) );
  XNOR2V0_8TH40 U1168 ( .A1(inst_i[12]), .A2(wb_cp0_waddr[1]), .ZN(n771) );
  CLKNV1_8TH40 U1169 ( .I(n231), .ZN(n1012) );
  AOI222V0_8TH40 U1170 ( .A1(df_memex_hi[0]), .A2(n259), .B1(df_wbex_hi[0]), 
        .B2(n260), .C1(hi_i[0]), .C2(n261), .ZN(n231) );
  I2NOR3V1_8TH40 U1171 ( .A1(df_wbex_hilo_we), .A2(n777), .B(df_memex_hilo_we), 
        .ZN(n260) );
  AND2V0_8TH40 U1172 ( .A1(df_memex_hilo_we), .A2(n777), .Z(n259) );
  CLKNV1_8TH40 U1173 ( .I(n257), .ZN(n289) );
  NAND4V0P5_8TH40 U1174 ( .A1(n757), .A2(n742), .A3(n234), .A4(n764), .ZN(n257) );
  NOR3V0P5_8TH40 U1175 ( .A1(n778), .A2(inst_class[2]), .A3(n763), .ZN(n757)
         );
  CLKNAND2V1_8TH40 U1176 ( .A1(n784), .A2(n236), .ZN(n346) );
  I2NOR3V1_8TH40 U1177 ( .A1(gpr1_data[5]), .A2(n395), .B(gpr1_data[4]), .ZN(
        n617) );
  CLKNV1_8TH40 U1178 ( .I(n458), .ZN(n397) );
  NAND3V0P5_8TH40 U1179 ( .A1(n786), .A2(n914), .A3(n395), .ZN(n458) );
  NOR2V0P5_8TH40 U1180 ( .A1(gpr1_data[24]), .A2(n1021), .ZN(n785) );
  OA221V0_8TH40 U1181 ( .A1(gpr1_data[16]), .A2(n350), .B1(gpr1_data[22]), 
        .B2(n386), .C(n787), .Z(n390) );
  AOAI211V0_8TH40 U1182 ( .A1(gpr1_data[19]), .A2(n1028), .B(n1026), .C(n618), 
        .ZN(n787) );
  AOAOAOI211111V0_8TH40 U1183 ( .A1(gpr1_data[27]), .A2(n1020), .B(n1018), .C(
        gpr1_data[29]), .D(n1016), .E(gpr1_data[31]), .F(n352), .ZN(n782) );
  AND3V0_8TH40 U1184 ( .A1(n786), .A2(n395), .A3(gpr1_data[2]), .Z(n325) );
  NOR3V0P5_8TH40 U1185 ( .A1(n1040), .A2(n1039), .A3(n388), .ZN(n395) );
  CLKNV1_8TH40 U1186 ( .I(n396), .ZN(n786) );
  NAND3V0P5_8TH40 U1187 ( .A1(gpr1_data[3]), .A2(gpr1_data[4]), .A3(
        gpr1_data[5]), .ZN(n396) );
  CLKNV1_8TH40 U1188 ( .I(n388), .ZN(n790) );
  NAND3V0P5_8TH40 U1189 ( .A1(n623), .A2(gpr1_data[10]), .A3(n348), .ZN(n388)
         );
  NOR2V0P5_8TH40 U1190 ( .A1(n1038), .A2(n1037), .ZN(n623) );
  AOAI211V0_8TH40 U1191 ( .A1(gpr1_data[9]), .A2(n1038), .B(n1036), .C(n348), 
        .ZN(n789) );
  CLKNV1_8TH40 U1192 ( .I(n622), .ZN(n348) );
  NAND3V0P5_8TH40 U1193 ( .A1(n464), .A2(gpr1_data[11]), .A3(n465), .ZN(n622)
         );
  CLKNV1_8TH40 U1194 ( .I(n626), .ZN(n465) );
  CLKNAND2V1_8TH40 U1195 ( .A1(n351), .A2(gpr1_data[14]), .ZN(n626) );
  NOR2V0P5_8TH40 U1196 ( .A1(n1034), .A2(n1033), .ZN(n464) );
  AOAI211V0_8TH40 U1197 ( .A1(gpr1_data[13]), .A2(n1034), .B(n1032), .C(n351), 
        .ZN(n788) );
  NOR3V0P5_8TH40 U1198 ( .A1(n1031), .A2(n1030), .A3(n350), .ZN(n351) );
  NAND3V0P5_8TH40 U1199 ( .A1(n624), .A2(gpr1_data[17]), .A3(n461), .ZN(n350)
         );
  INOR2V0_8TH40 U1200 ( .A1(n618), .B1(n1026), .ZN(n461) );
  NOR3V0P5_8TH40 U1201 ( .A1(n1025), .A2(n1024), .A3(n386), .ZN(n618) );
  CLKNAND2V1_8TH40 U1202 ( .A1(n383), .A2(gpr1_data[23]), .ZN(n386) );
  I2NOR3V1_8TH40 U1203 ( .A1(gpr1_data[24]), .A2(n625), .B(n1021), .ZN(n383)
         );
  NOR3V0P5_8TH40 U1204 ( .A1(n1020), .A2(n1019), .A3(n467), .ZN(n625) );
  INAND3V0_8TH40 U1205 ( .A1(n616), .B1(gpr1_data[30]), .B2(gpr1_data[31]), 
        .ZN(n467) );
  CLKNAND2V1_8TH40 U1206 ( .A1(gpr1_data[28]), .A2(gpr1_data[29]), .ZN(n616)
         );
  CLKNV1_8TH40 U1207 ( .I(n462), .ZN(n624) );
  CLKNAND2V1_8TH40 U1208 ( .A1(gpr1_data[18]), .A2(gpr1_data[19]), .ZN(n462)
         );
  CLKNAND2V1_8TH40 U1209 ( .A1(n688), .A2(n2), .ZN(n299) );
  CLKNV1_8TH40 U1210 ( .I(n539), .ZN(n276) );
  NOR2V0P5_8TH40 U1211 ( .A1(n353), .A2(N1873), .ZN(n539) );
  CLKNAND2V1_8TH40 U1212 ( .A1(n696), .A2(n912), .ZN(n353) );
  NOR2V0P5_8TH40 U1213 ( .A1(n1042), .A2(N1872), .ZN(n696) );
  OR2V0_8TH40 U1214 ( .A1(n793), .A2(n794), .Z(n791) );
  AOI211V0_8TH40 U1215 ( .A1(n611), .A2(gpr1_data[22]), .B(n374), .C(n361), 
        .ZN(n796) );
  OAOAI2111V0_8TH40 U1216 ( .A1(n1040), .A2(gpr1_data[7]), .B(n1038), .C(n609), 
        .D(n381), .ZN(n798) );
  NAND3V0P5_8TH40 U1217 ( .A1(gpr1_data[0]), .A2(n913), .A3(n327), .ZN(n381)
         );
  CLKNV1_8TH40 U1218 ( .I(n401), .ZN(n327) );
  NAND3V0P5_8TH40 U1219 ( .A1(n402), .A2(n914), .A3(n455), .ZN(n401) );
  OAOI211V0_8TH40 U1220 ( .A1(n1036), .A2(gpr1_data[11]), .B(n1034), .C(n610), 
        .ZN(n797) );
  OAI221V0_8TH40 U1221 ( .A1(n1030), .A2(n359), .B1(n1028), .B2(n376), .C(n598), .ZN(n374) );
  CLKNAND2V1_8TH40 U1222 ( .A1(n450), .A2(gpr1_data[20]), .ZN(n598) );
  NOR3V0P5_8TH40 U1223 ( .A1(gpr1_data[21]), .A2(gpr1_data[22]), .A3(n378), 
        .ZN(n450) );
  CLKNV1_8TH40 U1224 ( .I(n611), .ZN(n378) );
  AND3V0_8TH40 U1225 ( .A1(n607), .A2(n1021), .A3(gpr1_data[24]), .Z(n799) );
  NAND3V0P5_8TH40 U1226 ( .A1(n402), .A2(gpr1_data[2]), .A3(n455), .ZN(n400)
         );
  NOR3V0P5_8TH40 U1227 ( .A1(gpr1_data[4]), .A2(gpr1_data[5]), .A3(
        gpr1_data[3]), .ZN(n402) );
  NAND3V0P5_8TH40 U1228 ( .A1(gpr1_data[4]), .A2(n1041), .A3(n455), .ZN(n597)
         );
  CLKNV1_8TH40 U1229 ( .I(n403), .ZN(n455) );
  NAND3V0P5_8TH40 U1230 ( .A1(n1040), .A2(n1039), .A3(n382), .ZN(n403) );
  NOR2V0P5_8TH40 U1231 ( .A1(n609), .A2(gpr1_data[8]), .ZN(n382) );
  NAND3V0P5_8TH40 U1232 ( .A1(n606), .A2(n1037), .A3(n446), .ZN(n609) );
  NOR2V0P5_8TH40 U1233 ( .A1(n610), .A2(gpr1_data[12]), .ZN(n446) );
  NAND3V0P5_8TH40 U1234 ( .A1(n1033), .A2(n1032), .A3(n360), .ZN(n610) );
  NOR3V0P5_8TH40 U1235 ( .A1(gpr1_data[15]), .A2(gpr1_data[16]), .A3(n359), 
        .ZN(n360) );
  NAND3V0P5_8TH40 U1236 ( .A1(n1029), .A2(n1028), .A3(n448), .ZN(n359) );
  CLKNV1_8TH40 U1237 ( .I(n376), .ZN(n448) );
  NAND3V0P5_8TH40 U1238 ( .A1(n377), .A2(n1026), .A3(n611), .ZN(n376) );
  NOR2V0P5_8TH40 U1239 ( .A1(n379), .A2(gpr1_data[23]), .ZN(n611) );
  NAND3V0P5_8TH40 U1240 ( .A1(n1022), .A2(n1021), .A3(n607), .ZN(n379) );
  INOR3V0_8TH40 U1241 ( .A1(n451), .B1(n454), .B2(n452), .ZN(n607) );
  CLKNAND2V1_8TH40 U1242 ( .A1(n1019), .A2(n1020), .ZN(n452) );
  CLKNAND2V1_8TH40 U1243 ( .A1(n1016), .A2(n1015), .ZN(n454) );
  NOR2V0P5_8TH40 U1244 ( .A1(gpr1_data[29]), .A2(gpr1_data[28]), .ZN(n451) );
  NOR3V0P5_8TH40 U1245 ( .A1(gpr1_data[21]), .A2(gpr1_data[22]), .A3(
        gpr1_data[19]), .ZN(n377) );
  CLKNV1_8TH40 U1246 ( .I(n447), .ZN(n606) );
  CLKNAND2V1_8TH40 U1247 ( .A1(n1035), .A2(n1036), .ZN(n447) );
  CLKNV1_8TH40 U1248 ( .I(n358), .ZN(n326) );
  CLKNAND2V1_8TH40 U1249 ( .A1(n784), .A2(n742), .ZN(n358) );
  I2NOR4V0_8TH40 U1250 ( .A1(n234), .A2(inst_type[7]), .B1(n792), .B2(n747), 
        .ZN(n784) );
  NOR3V0P5_8TH40 U1251 ( .A1(n778), .A2(inst_class[0]), .A3(n800), .ZN(n245)
         );
  CLKNV1_8TH40 U1252 ( .I(n792), .ZN(n805) );
  NAND4V0P5_8TH40 U1253 ( .A1(inst_class[2]), .A2(n763), .A3(n778), .A4(n777), 
        .ZN(n792) );
  CLKNV1_8TH40 U1254 ( .I(inst_class[1]), .ZN(n778) );
  I2NOR4V0_8TH40 U1255 ( .A1(inst_type[4]), .A2(inst_type[6]), .B1(n806), .B2(
        n807), .ZN(n804) );
  OAI21V0_8TH40 U1256 ( .A1(n808), .A2(n809), .B(n664), .ZN(n252) );
  INAND3V0_8TH40 U1257 ( .A1(n809), .B1(inst_type[0]), .B2(inst_type[1]), .ZN(
        n664) );
  NAND4V0P5_8TH40 U1258 ( .A1(n743), .A2(n810), .A3(n758), .A4(n747), .ZN(n809) );
  NOR2V0P5_8TH40 U1259 ( .A1(rst), .A2(inst_type[7]), .ZN(n811) );
  NOR3V0P5_8TH40 U1260 ( .A1(n800), .A2(inst_class[1]), .A3(n763), .ZN(n251)
         );
  CLKNV1_8TH40 U1261 ( .I(inst_class[0]), .ZN(n763) );
  CLKNV1_8TH40 U1262 ( .I(inst_class[2]), .ZN(n800) );
  MUX2NV0_8TH40 U1263 ( .I0(n819), .I1(n807), .S(N1574), .ZN(n818) );
  CLKNAND2V1_8TH40 U1264 ( .A1(n742), .A2(n760), .ZN(n819) );
  CLKXOR2V2_8TH40 U1265 ( .A1(n793), .A2(inst_type[1]), .Z(n817) );
  MUX2NV0_8TH40 U1266 ( .I0(n822), .I1(N96), .S(inst_type[0]), .ZN(n793) );
  IOA22V0_8TH40 U1267 ( .B1(gpr2_data[31]), .B2(n1015), .A1(n823), .A2(
        sum_res[31]), .ZN(n822) );
  CKMUX2V2_8TH40 U1268 ( .I0(n742), .I1(n236), .S(N1574), .Z(n820) );
  CLKNAND2V1_8TH40 U1269 ( .A1(inst_type[6]), .A2(n235), .ZN(n812) );
  NOR2V0P5_8TH40 U1270 ( .A1(div_done), .A2(n18), .ZN(div_start) );
  NOR2V0P5_8TH40 U1271 ( .A1(n1064), .A2(n18), .ZN(div_opdata2[9]) );
  CLKNV1_8TH40 U1272 ( .I(gpr2_data[9]), .ZN(n1064) );
  NOR2V0P5_8TH40 U1273 ( .A1(n1065), .A2(n18), .ZN(div_opdata2[8]) );
  CLKNV1_8TH40 U1274 ( .I(gpr2_data[8]), .ZN(n1065) );
  NOR2V0P5_8TH40 U1275 ( .A1(n1066), .A2(n18), .ZN(div_opdata2[7]) );
  CLKNV1_8TH40 U1276 ( .I(gpr2_data[7]), .ZN(n1066) );
  NOR2V0P5_8TH40 U1277 ( .A1(n1067), .A2(n18), .ZN(div_opdata2[6]) );
  CLKNV1_8TH40 U1278 ( .I(gpr2_data[6]), .ZN(n1067) );
  NOR2V0P5_8TH40 U1279 ( .A1(n1068), .A2(n18), .ZN(div_opdata2[5]) );
  CLKNV1_8TH40 U1280 ( .I(gpr2_data[5]), .ZN(n1068) );
  NOR2V0P5_8TH40 U1281 ( .A1(n1069), .A2(n18), .ZN(div_opdata2[4]) );
  CLKNV1_8TH40 U1282 ( .I(gpr2_data[4]), .ZN(n1069) );
  NOR2V0P5_8TH40 U1283 ( .A1(n1070), .A2(n18), .ZN(div_opdata2[3]) );
  CLKNV1_8TH40 U1284 ( .I(gpr2_data[3]), .ZN(n1070) );
  NOR2V0P5_8TH40 U1285 ( .A1(n1042), .A2(n18), .ZN(div_opdata2[31]) );
  CLKNV1_8TH40 U1286 ( .I(gpr2_data[31]), .ZN(n1042) );
  NOR2V0P5_8TH40 U1287 ( .A1(n1043), .A2(n18), .ZN(div_opdata2[30]) );
  CLKNV1_8TH40 U1288 ( .I(gpr2_data[30]), .ZN(n1043) );
  NOR2V0P5_8TH40 U1289 ( .A1(n1071), .A2(n18), .ZN(div_opdata2[2]) );
  CLKNV1_8TH40 U1290 ( .I(gpr2_data[2]), .ZN(n1071) );
  NOR2V0P5_8TH40 U1291 ( .A1(n1044), .A2(n18), .ZN(div_opdata2[29]) );
  CLKNV1_8TH40 U1292 ( .I(gpr2_data[29]), .ZN(n1044) );
  NOR2V0P5_8TH40 U1293 ( .A1(n1045), .A2(n18), .ZN(div_opdata2[28]) );
  CLKNV1_8TH40 U1294 ( .I(gpr2_data[28]), .ZN(n1045) );
  NOR2V0P5_8TH40 U1295 ( .A1(n1046), .A2(n18), .ZN(div_opdata2[27]) );
  CLKNV1_8TH40 U1296 ( .I(gpr2_data[27]), .ZN(n1046) );
  NOR2V0P5_8TH40 U1297 ( .A1(n1047), .A2(n18), .ZN(div_opdata2[26]) );
  CLKNV1_8TH40 U1298 ( .I(gpr2_data[26]), .ZN(n1047) );
  NOR2V0P5_8TH40 U1299 ( .A1(n1048), .A2(n18), .ZN(div_opdata2[25]) );
  CLKNV1_8TH40 U1300 ( .I(gpr2_data[25]), .ZN(n1048) );
  NOR2V0P5_8TH40 U1301 ( .A1(n1049), .A2(n18), .ZN(div_opdata2[24]) );
  CLKNV1_8TH40 U1302 ( .I(gpr2_data[24]), .ZN(n1049) );
  NOR2V0P5_8TH40 U1303 ( .A1(n1050), .A2(n18), .ZN(div_opdata2[23]) );
  CLKNV1_8TH40 U1304 ( .I(gpr2_data[23]), .ZN(n1050) );
  NOR2V0P5_8TH40 U1305 ( .A1(n1051), .A2(n18), .ZN(div_opdata2[22]) );
  CLKNV1_8TH40 U1306 ( .I(gpr2_data[22]), .ZN(n1051) );
  NOR2V0P5_8TH40 U1307 ( .A1(n1052), .A2(n18), .ZN(div_opdata2[21]) );
  CLKNV1_8TH40 U1308 ( .I(gpr2_data[21]), .ZN(n1052) );
  NOR2V0P5_8TH40 U1309 ( .A1(n1053), .A2(n18), .ZN(div_opdata2[20]) );
  CLKNV1_8TH40 U1310 ( .I(gpr2_data[20]), .ZN(n1053) );
  NOR2V0P5_8TH40 U1311 ( .A1(n1072), .A2(n18), .ZN(div_opdata2[1]) );
  CLKNV1_8TH40 U1312 ( .I(gpr2_data[1]), .ZN(n1072) );
  NOR2V0P5_8TH40 U1313 ( .A1(n1054), .A2(n18), .ZN(div_opdata2[19]) );
  CLKNV1_8TH40 U1314 ( .I(gpr2_data[19]), .ZN(n1054) );
  NOR2V0P5_8TH40 U1315 ( .A1(n1055), .A2(n18), .ZN(div_opdata2[18]) );
  CLKNV1_8TH40 U1316 ( .I(gpr2_data[18]), .ZN(n1055) );
  NOR2V0P5_8TH40 U1317 ( .A1(n1056), .A2(n18), .ZN(div_opdata2[17]) );
  CLKNV1_8TH40 U1318 ( .I(gpr2_data[17]), .ZN(n1056) );
  NOR2V0P5_8TH40 U1319 ( .A1(n1057), .A2(n18), .ZN(div_opdata2[16]) );
  CLKNV1_8TH40 U1320 ( .I(gpr2_data[16]), .ZN(n1057) );
  NOR2V0P5_8TH40 U1321 ( .A1(n1058), .A2(n18), .ZN(div_opdata2[15]) );
  CLKNV1_8TH40 U1322 ( .I(gpr2_data[15]), .ZN(n1058) );
  NOR2V0P5_8TH40 U1323 ( .A1(n1059), .A2(n18), .ZN(div_opdata2[14]) );
  CLKNV1_8TH40 U1324 ( .I(gpr2_data[14]), .ZN(n1059) );
  NOR2V0P5_8TH40 U1325 ( .A1(n1060), .A2(n18), .ZN(div_opdata2[13]) );
  CLKNV1_8TH40 U1326 ( .I(gpr2_data[13]), .ZN(n1060) );
  NOR2V0P5_8TH40 U1327 ( .A1(n1061), .A2(n18), .ZN(div_opdata2[12]) );
  CLKNV1_8TH40 U1328 ( .I(gpr2_data[12]), .ZN(n1061) );
  NOR2V0P5_8TH40 U1329 ( .A1(n1062), .A2(n18), .ZN(div_opdata2[11]) );
  CLKNV1_8TH40 U1330 ( .I(gpr2_data[11]), .ZN(n1062) );
  NOR2V0P5_8TH40 U1331 ( .A1(n1063), .A2(n18), .ZN(div_opdata2[10]) );
  CLKNV1_8TH40 U1332 ( .I(gpr2_data[10]), .ZN(n1063) );
  NOR2V0P5_8TH40 U1333 ( .A1(n1073), .A2(n18), .ZN(div_opdata2[0]) );
  CLKNV1_8TH40 U1334 ( .I(gpr2_data[0]), .ZN(n1073) );
  NOR2V0P5_8TH40 U1335 ( .A1(n1037), .A2(n18), .ZN(div_opdata1[9]) );
  NOR2V0P5_8TH40 U1336 ( .A1(n1038), .A2(n18), .ZN(div_opdata1[8]) );
  NOR2V0P5_8TH40 U1337 ( .A1(n1039), .A2(n18), .ZN(div_opdata1[7]) );
  NOR2V0P5_8TH40 U1338 ( .A1(n1040), .A2(n18), .ZN(div_opdata1[6]) );
  NOR2V0P5_8TH40 U1339 ( .A1(n1041), .A2(n18), .ZN(div_opdata1[5]) );
  NOR2V0P5_8TH40 U1340 ( .A1(n916), .A2(n18), .ZN(div_opdata1[4]) );
  NOR2V0P5_8TH40 U1341 ( .A1(n915), .A2(n18), .ZN(div_opdata1[3]) );
  NOR2V0P5_8TH40 U1342 ( .A1(n1015), .A2(n18), .ZN(div_opdata1[31]) );
  NOR2V0P5_8TH40 U1343 ( .A1(n1016), .A2(n18), .ZN(div_opdata1[30]) );
  NOR2V0P5_8TH40 U1344 ( .A1(n914), .A2(n18), .ZN(div_opdata1[2]) );
  NOR2V0P5_8TH40 U1345 ( .A1(n1017), .A2(n18), .ZN(div_opdata1[29]) );
  NOR2V0P5_8TH40 U1346 ( .A1(n1018), .A2(n18), .ZN(div_opdata1[28]) );
  NOR2V0P5_8TH40 U1347 ( .A1(n1019), .A2(n18), .ZN(div_opdata1[27]) );
  NOR2V0P5_8TH40 U1348 ( .A1(n1020), .A2(n18), .ZN(div_opdata1[26]) );
  NOR2V0P5_8TH40 U1349 ( .A1(n1021), .A2(n18), .ZN(div_opdata1[25]) );
  NOR2V0P5_8TH40 U1350 ( .A1(n1022), .A2(n18), .ZN(div_opdata1[24]) );
  NOR2V0P5_8TH40 U1351 ( .A1(n1023), .A2(n18), .ZN(div_opdata1[23]) );
  NOR2V0P5_8TH40 U1352 ( .A1(n1024), .A2(n18), .ZN(div_opdata1[22]) );
  NOR2V0P5_8TH40 U1353 ( .A1(n1025), .A2(n18), .ZN(div_opdata1[21]) );
  NOR2V0P5_8TH40 U1354 ( .A1(n1026), .A2(n18), .ZN(div_opdata1[20]) );
  NOR2V0P5_8TH40 U1355 ( .A1(n913), .A2(n18), .ZN(div_opdata1[1]) );
  NOR2V0P5_8TH40 U1356 ( .A1(n1027), .A2(n18), .ZN(div_opdata1[19]) );
  NOR2V0P5_8TH40 U1357 ( .A1(n1028), .A2(n18), .ZN(div_opdata1[18]) );
  NOR2V0P5_8TH40 U1358 ( .A1(n1029), .A2(n18), .ZN(div_opdata1[17]) );
  NOR2V0P5_8TH40 U1359 ( .A1(n1030), .A2(n18), .ZN(div_opdata1[16]) );
  NOR2V0P5_8TH40 U1360 ( .A1(n1031), .A2(n18), .ZN(div_opdata1[15]) );
  NOR2V0P5_8TH40 U1361 ( .A1(n1032), .A2(n18), .ZN(div_opdata1[14]) );
  NOR2V0P5_8TH40 U1362 ( .A1(n1033), .A2(n18), .ZN(div_opdata1[13]) );
  NOR2V0P5_8TH40 U1363 ( .A1(n1034), .A2(n18), .ZN(div_opdata1[12]) );
  NOR2V0P5_8TH40 U1364 ( .A1(n1035), .A2(n18), .ZN(div_opdata1[11]) );
  NOR2V0P5_8TH40 U1365 ( .A1(n1036), .A2(n18), .ZN(div_opdata1[10]) );
  NOR2V0P5_8TH40 U1366 ( .A1(n912), .A2(n18), .ZN(div_opdata1[0]) );
  NAND3V0P5_8TH40 U1367 ( .A1(n235), .A2(n238), .A3(n759), .ZN(n18) );
  NOR2V0P5_8TH40 U1368 ( .A1(n806), .A2(rst), .ZN(n235) );
  NOR2V0P5_8TH40 U1369 ( .A1(n1037), .A2(n824), .ZN(cp0_wdata[9]) );
  CLKNV1_8TH40 U1370 ( .I(gpr1_data[9]), .ZN(n1037) );
  NOR2V0P5_8TH40 U1371 ( .A1(n1038), .A2(n824), .ZN(cp0_wdata[8]) );
  CLKNV1_8TH40 U1372 ( .I(gpr1_data[8]), .ZN(n1038) );
  NOR2V0P5_8TH40 U1373 ( .A1(n1039), .A2(n824), .ZN(cp0_wdata[7]) );
  CLKNV1_8TH40 U1374 ( .I(gpr1_data[7]), .ZN(n1039) );
  NOR2V0P5_8TH40 U1375 ( .A1(n1040), .A2(n824), .ZN(cp0_wdata[6]) );
  CLKNV1_8TH40 U1376 ( .I(gpr1_data[6]), .ZN(n1040) );
  NOR2V0P5_8TH40 U1377 ( .A1(n1041), .A2(n824), .ZN(cp0_wdata[5]) );
  CLKNV1_8TH40 U1378 ( .I(gpr1_data[5]), .ZN(n1041) );
  NOR2V0P5_8TH40 U1379 ( .A1(n916), .A2(n824), .ZN(cp0_wdata[4]) );
  CLKNV1_8TH40 U1380 ( .I(gpr1_data[4]), .ZN(n916) );
  NOR2V0P5_8TH40 U1381 ( .A1(n915), .A2(n824), .ZN(cp0_wdata[3]) );
  CLKNV1_8TH40 U1382 ( .I(gpr1_data[3]), .ZN(n915) );
  NOR2V0P5_8TH40 U1383 ( .A1(n1015), .A2(n824), .ZN(cp0_wdata[31]) );
  NOR2V0P5_8TH40 U1384 ( .A1(n1016), .A2(n824), .ZN(cp0_wdata[30]) );
  CLKNV1_8TH40 U1385 ( .I(gpr1_data[30]), .ZN(n1016) );
  NOR2V0P5_8TH40 U1386 ( .A1(n914), .A2(n824), .ZN(cp0_wdata[2]) );
  CLKNV1_8TH40 U1387 ( .I(gpr1_data[2]), .ZN(n914) );
  NOR2V0P5_8TH40 U1388 ( .A1(n1017), .A2(n824), .ZN(cp0_wdata[29]) );
  CLKNV1_8TH40 U1389 ( .I(gpr1_data[29]), .ZN(n1017) );
  NOR2V0P5_8TH40 U1390 ( .A1(n1018), .A2(n824), .ZN(cp0_wdata[28]) );
  CLKNV1_8TH40 U1391 ( .I(gpr1_data[28]), .ZN(n1018) );
  NOR2V0P5_8TH40 U1392 ( .A1(n1019), .A2(n824), .ZN(cp0_wdata[27]) );
  CLKNV1_8TH40 U1393 ( .I(gpr1_data[27]), .ZN(n1019) );
  NOR2V0P5_8TH40 U1394 ( .A1(n1020), .A2(n824), .ZN(cp0_wdata[26]) );
  CLKNV1_8TH40 U1395 ( .I(gpr1_data[26]), .ZN(n1020) );
  NOR2V0P5_8TH40 U1396 ( .A1(n1021), .A2(n824), .ZN(cp0_wdata[25]) );
  CLKNV1_8TH40 U1397 ( .I(gpr1_data[25]), .ZN(n1021) );
  NOR2V0P5_8TH40 U1398 ( .A1(n1022), .A2(n824), .ZN(cp0_wdata[24]) );
  CLKNV1_8TH40 U1399 ( .I(gpr1_data[24]), .ZN(n1022) );
  NOR2V0P5_8TH40 U1400 ( .A1(n1023), .A2(n824), .ZN(cp0_wdata[23]) );
  CLKNV1_8TH40 U1401 ( .I(gpr1_data[23]), .ZN(n1023) );
  NOR2V0P5_8TH40 U1402 ( .A1(n1024), .A2(n824), .ZN(cp0_wdata[22]) );
  CLKNV1_8TH40 U1403 ( .I(gpr1_data[22]), .ZN(n1024) );
  NOR2V0P5_8TH40 U1404 ( .A1(n1025), .A2(n824), .ZN(cp0_wdata[21]) );
  CLKNV1_8TH40 U1405 ( .I(gpr1_data[21]), .ZN(n1025) );
  NOR2V0P5_8TH40 U1406 ( .A1(n1026), .A2(n824), .ZN(cp0_wdata[20]) );
  CLKNV1_8TH40 U1407 ( .I(gpr1_data[20]), .ZN(n1026) );
  NOR2V0P5_8TH40 U1408 ( .A1(n913), .A2(n824), .ZN(cp0_wdata[1]) );
  CLKNV1_8TH40 U1409 ( .I(gpr1_data[1]), .ZN(n913) );
  NOR2V0P5_8TH40 U1410 ( .A1(n1027), .A2(n824), .ZN(cp0_wdata[19]) );
  CLKNV1_8TH40 U1411 ( .I(gpr1_data[19]), .ZN(n1027) );
  NOR2V0P5_8TH40 U1412 ( .A1(n1028), .A2(n824), .ZN(cp0_wdata[18]) );
  CLKNV1_8TH40 U1413 ( .I(gpr1_data[18]), .ZN(n1028) );
  NOR2V0P5_8TH40 U1414 ( .A1(n1029), .A2(n824), .ZN(cp0_wdata[17]) );
  CLKNV1_8TH40 U1415 ( .I(gpr1_data[17]), .ZN(n1029) );
  NOR2V0P5_8TH40 U1416 ( .A1(n1030), .A2(n824), .ZN(cp0_wdata[16]) );
  CLKNV1_8TH40 U1417 ( .I(gpr1_data[16]), .ZN(n1030) );
  NOR2V0P5_8TH40 U1418 ( .A1(n1031), .A2(n824), .ZN(cp0_wdata[15]) );
  CLKNV1_8TH40 U1419 ( .I(gpr1_data[15]), .ZN(n1031) );
  NOR2V0P5_8TH40 U1420 ( .A1(n1032), .A2(n824), .ZN(cp0_wdata[14]) );
  CLKNV1_8TH40 U1421 ( .I(gpr1_data[14]), .ZN(n1032) );
  NOR2V0P5_8TH40 U1422 ( .A1(n1033), .A2(n824), .ZN(cp0_wdata[13]) );
  CLKNV1_8TH40 U1423 ( .I(gpr1_data[13]), .ZN(n1033) );
  NOR2V0P5_8TH40 U1424 ( .A1(n1034), .A2(n824), .ZN(cp0_wdata[12]) );
  CLKNV1_8TH40 U1425 ( .I(gpr1_data[12]), .ZN(n1034) );
  NOR2V0P5_8TH40 U1426 ( .A1(n1035), .A2(n824), .ZN(cp0_wdata[11]) );
  CLKNV1_8TH40 U1427 ( .I(gpr1_data[11]), .ZN(n1035) );
  NOR2V0P5_8TH40 U1428 ( .A1(n1036), .A2(n824), .ZN(cp0_wdata[10]) );
  CLKNV1_8TH40 U1429 ( .I(gpr1_data[10]), .ZN(n1036) );
  NOR2V0P5_8TH40 U1430 ( .A1(n912), .A2(n824), .ZN(cp0_wdata[0]) );
  CLKNV1_8TH40 U1431 ( .I(gpr1_data[0]), .ZN(n912) );
  AND2V0_8TH40 U1432 ( .A1(inst_i[15]), .A2(cp0_we), .Z(cp0_waddr[4]) );
  AND2V0_8TH40 U1433 ( .A1(inst_i[14]), .A2(cp0_we), .Z(cp0_waddr[3]) );
  AND2V0_8TH40 U1434 ( .A1(inst_i[13]), .A2(cp0_we), .Z(cp0_waddr[2]) );
  CLKNV1_8TH40 U1435 ( .I(n824), .ZN(cp0_we) );
  INOR2V0_8TH40 U1436 ( .A1(inst_i[12]), .B1(n824), .ZN(cp0_waddr[1]) );
  INOR2V0_8TH40 U1437 ( .A1(inst_i[11]), .B1(n824), .ZN(cp0_waddr[0]) );
  NOR3V0P5_8TH40 U1438 ( .A1(n816), .A2(rst), .A3(inst_type[4]), .ZN(n825) );
  CLKNV1_8TH40 U1439 ( .I(n826), .ZN(n816) );
  CKMUX2V2_8TH40 U1440 ( .I0(N69), .I1(gpr2_data[9]), .S(n827), .Z(
        com_gpr2_data[9]) );
  CKMUX2V2_8TH40 U1441 ( .I0(N68), .I1(gpr2_data[8]), .S(n827), .Z(
        com_gpr2_data[8]) );
  CKMUX2V2_8TH40 U1442 ( .I0(N67), .I1(gpr2_data[7]), .S(n827), .Z(
        com_gpr2_data[7]) );
  CKMUX2V2_8TH40 U1443 ( .I0(N66), .I1(gpr2_data[6]), .S(n827), .Z(
        com_gpr2_data[6]) );
  CKMUX2V2_8TH40 U1444 ( .I0(N65), .I1(gpr2_data[5]), .S(n827), .Z(
        com_gpr2_data[5]) );
  CKMUX2V2_8TH40 U1445 ( .I0(N64), .I1(gpr2_data[4]), .S(n827), .Z(
        com_gpr2_data[4]) );
  CKMUX2V2_8TH40 U1446 ( .I0(N63), .I1(gpr2_data[3]), .S(n827), .Z(
        com_gpr2_data[3]) );
  CKMUX2V2_8TH40 U1447 ( .I0(N90), .I1(gpr2_data[30]), .S(n827), .Z(
        com_gpr2_data[30]) );
  CKMUX2V2_8TH40 U1448 ( .I0(N62), .I1(gpr2_data[2]), .S(n827), .Z(
        com_gpr2_data[2]) );
  CKMUX2V2_8TH40 U1449 ( .I0(N89), .I1(gpr2_data[29]), .S(n827), .Z(
        com_gpr2_data[29]) );
  CKMUX2V2_8TH40 U1450 ( .I0(N88), .I1(gpr2_data[28]), .S(n827), .Z(
        com_gpr2_data[28]) );
  CKMUX2V2_8TH40 U1451 ( .I0(N87), .I1(gpr2_data[27]), .S(n827), .Z(
        com_gpr2_data[27]) );
  CKMUX2V2_8TH40 U1452 ( .I0(N86), .I1(gpr2_data[26]), .S(n827), .Z(
        com_gpr2_data[26]) );
  CKMUX2V2_8TH40 U1453 ( .I0(N85), .I1(gpr2_data[25]), .S(n827), .Z(
        com_gpr2_data[25]) );
  CKMUX2V2_8TH40 U1454 ( .I0(N84), .I1(gpr2_data[24]), .S(n827), .Z(
        com_gpr2_data[24]) );
  CKMUX2V2_8TH40 U1455 ( .I0(N83), .I1(gpr2_data[23]), .S(n827), .Z(
        com_gpr2_data[23]) );
  CKMUX2V2_8TH40 U1456 ( .I0(N82), .I1(gpr2_data[22]), .S(n827), .Z(
        com_gpr2_data[22]) );
  CKMUX2V2_8TH40 U1457 ( .I0(N81), .I1(gpr2_data[21]), .S(n827), .Z(
        com_gpr2_data[21]) );
  CKMUX2V2_8TH40 U1458 ( .I0(N80), .I1(gpr2_data[20]), .S(n827), .Z(
        com_gpr2_data[20]) );
  CKMUX2V2_8TH40 U1459 ( .I0(N61), .I1(gpr2_data[1]), .S(n827), .Z(
        com_gpr2_data[1]) );
  CKMUX2V2_8TH40 U1460 ( .I0(N79), .I1(gpr2_data[19]), .S(n827), .Z(
        com_gpr2_data[19]) );
  CKMUX2V2_8TH40 U1461 ( .I0(N78), .I1(gpr2_data[18]), .S(n827), .Z(
        com_gpr2_data[18]) );
  CKMUX2V2_8TH40 U1462 ( .I0(N77), .I1(gpr2_data[17]), .S(n827), .Z(
        com_gpr2_data[17]) );
  CKMUX2V2_8TH40 U1463 ( .I0(N76), .I1(gpr2_data[16]), .S(n827), .Z(
        com_gpr2_data[16]) );
  CKMUX2V2_8TH40 U1464 ( .I0(N75), .I1(gpr2_data[15]), .S(n827), .Z(
        com_gpr2_data[15]) );
  CKMUX2V2_8TH40 U1465 ( .I0(N74), .I1(gpr2_data[14]), .S(n827), .Z(
        com_gpr2_data[14]) );
  CKMUX2V2_8TH40 U1466 ( .I0(N73), .I1(gpr2_data[13]), .S(n827), .Z(
        com_gpr2_data[13]) );
  CKMUX2V2_8TH40 U1467 ( .I0(N72), .I1(gpr2_data[12]), .S(n827), .Z(
        com_gpr2_data[12]) );
  CKMUX2V2_8TH40 U1468 ( .I0(N71), .I1(gpr2_data[11]), .S(n827), .Z(
        com_gpr2_data[11]) );
  CKMUX2V2_8TH40 U1469 ( .I0(N70), .I1(gpr2_data[10]), .S(n827), .Z(
        com_gpr2_data[10]) );
  AOAI211V0_8TH40 U1470 ( .A1(n830), .A2(n802), .B(n803), .C(n745), .ZN(n829)
         );
  CLKNV1_8TH40 U1471 ( .I(n831), .ZN(n803) );
  INAND2V0_8TH40 U1472 ( .A1(sum_res[31]), .B1(n917), .ZN(n833) );
  CLKNV1_8TH40 U1473 ( .I(n834), .ZN(n917) );
  CLKNAND2V1_8TH40 U1474 ( .A1(sum_res[31]), .A2(n834), .ZN(n832) );
  MUX2NV0_8TH40 U1475 ( .I0(N91), .I1(gpr2_data[31]), .S(n827), .ZN(n834) );
  I2NOR4V0_8TH40 U1476 ( .A1(n760), .A2(inst_type[6]), .B1(inst_type[4]), .B2(
        n806), .ZN(n836) );
  INOR2V0_8TH40 U1477 ( .A1(n810), .B1(n815), .ZN(n234) );
  CLKNV1_8TH40 U1478 ( .I(n238), .ZN(n815) );
  NOR2V0P5_8TH40 U1479 ( .A1(inst_type[2]), .A2(inst_type[3]), .ZN(n810) );
  NOR2V0P5_8TH40 U1480 ( .A1(n762), .A2(inst_type[2]), .ZN(n802) );
  CLKNAND2V1_8TH40 U1481 ( .A1(n826), .A2(n758), .ZN(n762) );
  NOR2V0P5_8TH40 U1482 ( .A1(n747), .A2(inst_type[7]), .ZN(n826) );
  CLKNV1_8TH40 U1483 ( .I(inst_type[5]), .ZN(n747) );
  NOR3V0P5_8TH40 U1484 ( .A1(n745), .A2(rst), .A3(n831), .ZN(N2186) );
  NOR2V0P5_8TH40 U1485 ( .A1(n806), .A2(n746), .ZN(n837) );
  CLKNV1_8TH40 U1486 ( .I(n764), .ZN(n806) );
  CLKNV1_8TH40 U1487 ( .I(inst_type[3]), .ZN(n745) );
  INAND2V0_8TH40 U1488 ( .A1(N1412), .B1(n838), .ZN(N1416) );
  I2NOR3V1_8TH40 U1489 ( .A1(n3), .A2(cycl_cnt_i[0]), .B(cycl_cnt_i[1]), .ZN(
        N1412) );
  AOI22V0_8TH40 U1490 ( .A1(mul_res_tmp[63]), .A2(n843), .B1(N666), .B2(n844), 
        .ZN(n149) );
  AOI22V0_8TH40 U1491 ( .A1(mul_res_tmp[43]), .A2(n843), .B1(N646), .B2(n844), 
        .ZN(n227) );
  AOI22V0_8TH40 U1492 ( .A1(mul_res_tmp[42]), .A2(n843), .B1(N645), .B2(n844), 
        .ZN(n230) );
  AOI22V0_8TH40 U1493 ( .A1(mul_res_tmp[41]), .A2(n843), .B1(N644), .B2(n844), 
        .ZN(n124) );
  AOI22V0_8TH40 U1494 ( .A1(mul_res_tmp[40]), .A2(n843), .B1(N643), .B2(n844), 
        .ZN(n127) );
  AOI22V0_8TH40 U1495 ( .A1(mul_res_tmp[39]), .A2(n843), .B1(N642), .B2(n844), 
        .ZN(n131) );
  AOI22V0_8TH40 U1496 ( .A1(mul_res_tmp[38]), .A2(n843), .B1(N641), .B2(n844), 
        .ZN(n134) );
  AOI22V0_8TH40 U1497 ( .A1(mul_res_tmp[37]), .A2(n843), .B1(N640), .B2(n844), 
        .ZN(n138) );
  AOI22V0_8TH40 U1498 ( .A1(mul_res_tmp[36]), .A2(n843), .B1(N639), .B2(n844), 
        .ZN(n141) );
  AOI22V0_8TH40 U1499 ( .A1(mul_res_tmp[35]), .A2(n843), .B1(N638), .B2(n844), 
        .ZN(n145) );
  AOI22V0_8TH40 U1500 ( .A1(mul_res_tmp[34]), .A2(n843), .B1(N637), .B2(n844), 
        .ZN(n155) );
  AOI22V0_8TH40 U1501 ( .A1(mul_res_tmp[33]), .A2(n843), .B1(N636), .B2(n844), 
        .ZN(n196) );
  AOI22V0_8TH40 U1502 ( .A1(mul_res_tmp[32]), .A2(n843), .B1(N635), .B2(n844), 
        .ZN(n237) );
  AOI22V0_8TH40 U1503 ( .A1(mul_res_tmp[31]), .A2(n843), .B1(N634), .B2(n844), 
        .ZN(n417) );
  AOI22V0_8TH40 U1504 ( .A1(mul_res_tmp[30]), .A2(n843), .B1(N633), .B2(n844), 
        .ZN(n425) );
  AOI22V0_8TH40 U1505 ( .A1(mul_res_tmp[23]), .A2(n843), .B1(N626), .B2(n844), 
        .ZN(n546) );
  AOI22V0_8TH40 U1506 ( .A1(mul_res_tmp[19]), .A2(n843), .B1(N622), .B2(n844), 
        .ZN(n633) );
  AOI22V0_8TH40 U1507 ( .A1(mul_res_tmp[18]), .A2(n843), .B1(N621), .B2(n844), 
        .ZN(n644) );
  AOI22V0_8TH40 U1508 ( .A1(mul_res_tmp[17]), .A2(n843), .B1(N620), .B2(n844), 
        .ZN(n654) );
  AOI22V0_8TH40 U1509 ( .A1(mul_res_tmp[16]), .A2(n843), .B1(N619), .B2(n844), 
        .ZN(n665) );
  AOI22V0_8TH40 U1510 ( .A1(mul_res_tmp[11]), .A2(n843), .B1(N614), .B2(n844), 
        .ZN(n717) );
  AOI22V0_8TH40 U1511 ( .A1(mul_res_tmp[3]), .A2(n843), .B1(N606), .B2(n844), 
        .ZN(n391) );
  AOI22V0_8TH40 U1512 ( .A1(mul_res_tmp[2]), .A2(n843), .B1(N605), .B2(n844), 
        .ZN(n468) );
  AOI22V0_8TH40 U1513 ( .A1(mul_res_tmp[1]), .A2(n843), .B1(N604), .B2(n844), 
        .ZN(n627) );
  AND2V0_8TH40 U1514 ( .A1(N1414), .A2(n1013), .Z(N1348) );
  AO22V0_8TH40 U1515 ( .A1(mul_res_tmp[0]), .A2(n843), .B1(N603), .B2(n844), 
        .Z(n1013) );
  I2NOR3V1_8TH40 U1516 ( .A1(n414), .A2(n35), .B(rst), .ZN(n844) );
  OAI21V0_8TH40 U1517 ( .A1(gpr2_data[31]), .A2(n1015), .B(n823), .ZN(n414) );
  CLKNAND2V1_8TH40 U1518 ( .A1(gpr2_data[31]), .A2(n1015), .ZN(n823) );
  CLKNV1_8TH40 U1519 ( .I(gpr1_data[31]), .ZN(n1015) );
  IAO21V0_8TH40 U1520 ( .A1(n755), .A2(n236), .B(n840), .ZN(n908) );
  NOR2V0P5_8TH40 U1521 ( .A1(n830), .A2(inst_type[1]), .ZN(n236) );
  NOR2V0P5_8TH40 U1522 ( .A1(inst_type[5]), .A2(inst_type[7]), .ZN(n764) );
  NOR2V0P5_8TH40 U1523 ( .A1(n746), .A2(inst_type[6]), .ZN(n238) );
  CLKNV1_8TH40 U1524 ( .I(inst_type[4]), .ZN(n746) );
  CLKNAND2V1_8TH40 U1525 ( .A1(n838), .A2(n842), .ZN(N1414) );
  NOR3V0P5_8TH40 U1526 ( .A1(cycl_cnt_i[0]), .A2(rst), .A3(cycl_cnt_i[1]), 
        .ZN(n909) );
  CLKNV1_8TH40 U1527 ( .I(rst), .ZN(n777) );
  NAND3V0P5_8TH40 U1528 ( .A1(n758), .A2(inst_type[5]), .A3(inst_type[7]), 
        .ZN(n840) );
  NOR2V0P5_8TH40 U1529 ( .A1(inst_type[4]), .A2(inst_type[6]), .ZN(n758) );
  CLKNV1_8TH40 U1530 ( .I(n794), .ZN(n759) );
  CLKNAND2V1_8TH40 U1531 ( .A1(inst_type[1]), .A2(n821), .ZN(n794) );
  NOR2V0P5_8TH40 U1532 ( .A1(cycl_cnt_i[1]), .A2(n839), .ZN(n910) );
  IAOI21V1_8TH40 U1533 ( .B1(n821), .B2(n742), .A(n807), .ZN(n839) );
  CLKNAND2V1_8TH40 U1534 ( .A1(n755), .A2(n760), .ZN(n807) );
  NOR2V0P5_8TH40 U1535 ( .A1(n748), .A2(inst_type[3]), .ZN(n760) );
  CLKNV1_8TH40 U1536 ( .I(n808), .ZN(n755) );
  CLKNAND2V1_8TH40 U1537 ( .A1(inst_type[1]), .A2(n830), .ZN(n808) );
  CLKNV1_8TH40 U1538 ( .I(inst_type[0]), .ZN(n830) );
  NOR2V0P5_8TH40 U1539 ( .A1(inst_type[0]), .A2(inst_type[1]), .ZN(n742) );
  CLKNV1_8TH40 U1540 ( .I(n239), .ZN(n821) );
  CLKNAND2V1_8TH40 U1541 ( .A1(inst_type[3]), .A2(n748), .ZN(n239) );
  CLKNV1_8TH40 U1542 ( .I(inst_type[2]), .ZN(n748) );
endmodule


module pipe_reg_exmem ( clk, rst, stall_ctrl, ex_gpr_we, ex_target_gpr, 
        ex_exe_result, ex_hi, ex_lo, ex_hilo_we, ex_hilo_tmp_i, ex_cycl_cnt_i, 
        ex_inst_type, ex_dmem_addr, ex_ls_data_tmp, ex_cp0_we, ex_cp0_waddr, 
        ex_cp0_wdata, ex_except_type, ex_cur_inst_addr, ex_inst_delayslot, 
        ex_hilo_tmp_o, ex_cycl_cnt_o, mem_gpr_we, mem_target_gpr, 
        mem_exe_result, mem_hi, mem_lo, mem_hilo_we, mem_inst_type, 
        mem_dmem_addr, mem_ls_data_tmp, mem_cp0_we, mem_cp0_waddr, 
        mem_cp0_wdata, mem_except_type, mem_cur_inst_addr, mem_inst_delayslot, 
        flush_BAR );
  input [5:0] stall_ctrl;
  input [4:0] ex_target_gpr;
  input [31:0] ex_exe_result;
  input [31:0] ex_hi;
  input [31:0] ex_lo;
  input [63:0] ex_hilo_tmp_i;
  input [1:0] ex_cycl_cnt_i;
  input [7:0] ex_inst_type;
  input [31:0] ex_dmem_addr;
  input [31:0] ex_ls_data_tmp;
  input [4:0] ex_cp0_waddr;
  input [31:0] ex_cp0_wdata;
  input [31:0] ex_except_type;
  input [31:0] ex_cur_inst_addr;
  output [63:0] ex_hilo_tmp_o;
  output [1:0] ex_cycl_cnt_o;
  output [4:0] mem_target_gpr;
  output [31:0] mem_exe_result;
  output [31:0] mem_hi;
  output [31:0] mem_lo;
  output [7:0] mem_inst_type;
  output [31:0] mem_dmem_addr;
  output [31:0] mem_ls_data_tmp;
  output [4:0] mem_cp0_waddr;
  output [31:0] mem_cp0_wdata;
  output [31:0] mem_except_type;
  output [31:0] mem_cur_inst_addr;
  input clk, rst, ex_gpr_we, ex_hilo_we, ex_cp0_we, ex_inst_delayslot,
         flush_BAR;
  output mem_gpr_we, mem_hilo_we, mem_cp0_we, mem_inst_delayslot;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n227, n228, n229, n230, n231,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n1, n2,
         n3, n4, n219, n220, n221, n222, n223, n224, n225, n226, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313;

  DQV4_8TH40 mem_cur_inst_addr_reg_31_ ( .D(n282), .CK(clk), .Q(
        mem_cur_inst_addr[31]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_30_ ( .D(n281), .CK(clk), .Q(
        mem_cur_inst_addr[30]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_29_ ( .D(n280), .CK(clk), .Q(
        mem_cur_inst_addr[29]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_28_ ( .D(n279), .CK(clk), .Q(
        mem_cur_inst_addr[28]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_27_ ( .D(n278), .CK(clk), .Q(
        mem_cur_inst_addr[27]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_26_ ( .D(n277), .CK(clk), .Q(
        mem_cur_inst_addr[26]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_25_ ( .D(n276), .CK(clk), .Q(
        mem_cur_inst_addr[25]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_24_ ( .D(n275), .CK(clk), .Q(
        mem_cur_inst_addr[24]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_23_ ( .D(n274), .CK(clk), .Q(
        mem_cur_inst_addr[23]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_22_ ( .D(n273), .CK(clk), .Q(
        mem_cur_inst_addr[22]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_21_ ( .D(n272), .CK(clk), .Q(
        mem_cur_inst_addr[21]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_20_ ( .D(n271), .CK(clk), .Q(
        mem_cur_inst_addr[20]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_19_ ( .D(n270), .CK(clk), .Q(
        mem_cur_inst_addr[19]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_18_ ( .D(n269), .CK(clk), .Q(
        mem_cur_inst_addr[18]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_17_ ( .D(n268), .CK(clk), .Q(
        mem_cur_inst_addr[17]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_16_ ( .D(n267), .CK(clk), .Q(
        mem_cur_inst_addr[16]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_15_ ( .D(n266), .CK(clk), .Q(
        mem_cur_inst_addr[15]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_14_ ( .D(n265), .CK(clk), .Q(
        mem_cur_inst_addr[14]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_13_ ( .D(n264), .CK(clk), .Q(
        mem_cur_inst_addr[13]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_12_ ( .D(n263), .CK(clk), .Q(
        mem_cur_inst_addr[12]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_11_ ( .D(n262), .CK(clk), .Q(
        mem_cur_inst_addr[11]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_10_ ( .D(n261), .CK(clk), .Q(
        mem_cur_inst_addr[10]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_9_ ( .D(n260), .CK(clk), .Q(
        mem_cur_inst_addr[9]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_8_ ( .D(n259), .CK(clk), .Q(
        mem_cur_inst_addr[8]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_7_ ( .D(n258), .CK(clk), .Q(
        mem_cur_inst_addr[7]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_6_ ( .D(n257), .CK(clk), .Q(
        mem_cur_inst_addr[6]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_5_ ( .D(n256), .CK(clk), .Q(
        mem_cur_inst_addr[5]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_4_ ( .D(n255), .CK(clk), .Q(
        mem_cur_inst_addr[4]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_3_ ( .D(n254), .CK(clk), .Q(
        mem_cur_inst_addr[3]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_2_ ( .D(n253), .CK(clk), .Q(
        mem_cur_inst_addr[2]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_1_ ( .D(n252), .CK(clk), .Q(
        mem_cur_inst_addr[1]) );
  DQV4_8TH40 mem_cur_inst_addr_reg_0_ ( .D(n251), .CK(clk), .Q(
        mem_cur_inst_addr[0]) );
  DQV4_8TH40 mem_except_type_reg_12_ ( .D(n231), .CK(clk), .Q(
        mem_except_type[12]) );
  DQV4_8TH40 mem_except_type_reg_11_ ( .D(n230), .CK(clk), .Q(
        mem_except_type[11]) );
  DQV4_8TH40 mem_except_type_reg_10_ ( .D(n229), .CK(clk), .Q(
        mem_except_type[10]) );
  DQV4_8TH40 mem_except_type_reg_9_ ( .D(n228), .CK(clk), .Q(
        mem_except_type[9]) );
  DQV4_8TH40 mem_except_type_reg_8_ ( .D(n227), .CK(clk), .Q(
        mem_except_type[8]) );
  DQV4_8TH40 mem_cp0_waddr_reg_4_ ( .D(n218), .CK(clk), .Q(mem_cp0_waddr[4])
         );
  DQV4_8TH40 mem_cp0_waddr_reg_3_ ( .D(n217), .CK(clk), .Q(mem_cp0_waddr[3])
         );
  DQV4_8TH40 mem_cp0_waddr_reg_2_ ( .D(n216), .CK(clk), .Q(mem_cp0_waddr[2])
         );
  DQV4_8TH40 mem_cp0_waddr_reg_1_ ( .D(n215), .CK(clk), .Q(mem_cp0_waddr[1])
         );
  DQV4_8TH40 mem_cp0_waddr_reg_0_ ( .D(n214), .CK(clk), .Q(mem_cp0_waddr[0])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_31_ ( .D(n213), .CK(clk), .Q(mem_cp0_wdata[31])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_30_ ( .D(n212), .CK(clk), .Q(mem_cp0_wdata[30])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_29_ ( .D(n211), .CK(clk), .Q(mem_cp0_wdata[29])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_28_ ( .D(n210), .CK(clk), .Q(mem_cp0_wdata[28])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_27_ ( .D(n209), .CK(clk), .Q(mem_cp0_wdata[27])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_26_ ( .D(n208), .CK(clk), .Q(mem_cp0_wdata[26])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_25_ ( .D(n207), .CK(clk), .Q(mem_cp0_wdata[25])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_24_ ( .D(n206), .CK(clk), .Q(mem_cp0_wdata[24])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_23_ ( .D(n205), .CK(clk), .Q(mem_cp0_wdata[23])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_22_ ( .D(n204), .CK(clk), .Q(mem_cp0_wdata[22])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_21_ ( .D(n203), .CK(clk), .Q(mem_cp0_wdata[21])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_20_ ( .D(n202), .CK(clk), .Q(mem_cp0_wdata[20])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_19_ ( .D(n201), .CK(clk), .Q(mem_cp0_wdata[19])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_18_ ( .D(n200), .CK(clk), .Q(mem_cp0_wdata[18])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_17_ ( .D(n199), .CK(clk), .Q(mem_cp0_wdata[17])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_16_ ( .D(n198), .CK(clk), .Q(mem_cp0_wdata[16])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_15_ ( .D(n197), .CK(clk), .Q(mem_cp0_wdata[15])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_14_ ( .D(n196), .CK(clk), .Q(mem_cp0_wdata[14])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_13_ ( .D(n195), .CK(clk), .Q(mem_cp0_wdata[13])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_12_ ( .D(n194), .CK(clk), .Q(mem_cp0_wdata[12])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_11_ ( .D(n193), .CK(clk), .Q(mem_cp0_wdata[11])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_10_ ( .D(n192), .CK(clk), .Q(mem_cp0_wdata[10])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_9_ ( .D(n191), .CK(clk), .Q(mem_cp0_wdata[9])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_8_ ( .D(n190), .CK(clk), .Q(mem_cp0_wdata[8])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_7_ ( .D(n189), .CK(clk), .Q(mem_cp0_wdata[7])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_6_ ( .D(n188), .CK(clk), .Q(mem_cp0_wdata[6])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_5_ ( .D(n187), .CK(clk), .Q(mem_cp0_wdata[5])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_4_ ( .D(n186), .CK(clk), .Q(mem_cp0_wdata[4])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_3_ ( .D(n185), .CK(clk), .Q(mem_cp0_wdata[3])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_2_ ( .D(n184), .CK(clk), .Q(mem_cp0_wdata[2])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_1_ ( .D(n183), .CK(clk), .Q(mem_cp0_wdata[1])
         );
  DQV4_8TH40 mem_cp0_wdata_reg_0_ ( .D(n182), .CK(clk), .Q(mem_cp0_wdata[0])
         );
  DQV4_8TH40 mem_inst_delayslot_reg ( .D(n181), .CK(clk), .Q(
        mem_inst_delayslot) );
  DQV4_8TH40 mem_gpr_we_reg ( .D(n180), .CK(clk), .Q(mem_gpr_we) );
  DQV4_8TH40 mem_target_gpr_reg_4_ ( .D(n179), .CK(clk), .Q(mem_target_gpr[4])
         );
  DQV4_8TH40 mem_target_gpr_reg_3_ ( .D(n178), .CK(clk), .Q(mem_target_gpr[3])
         );
  DQV4_8TH40 mem_target_gpr_reg_2_ ( .D(n177), .CK(clk), .Q(mem_target_gpr[2])
         );
  DQV4_8TH40 mem_target_gpr_reg_1_ ( .D(n176), .CK(clk), .Q(mem_target_gpr[1])
         );
  DQV4_8TH40 mem_target_gpr_reg_0_ ( .D(n175), .CK(clk), .Q(mem_target_gpr[0])
         );
  DQV4_8TH40 mem_exe_result_reg_31_ ( .D(n174), .CK(clk), .Q(
        mem_exe_result[31]) );
  DQV4_8TH40 mem_exe_result_reg_30_ ( .D(n173), .CK(clk), .Q(
        mem_exe_result[30]) );
  DQV4_8TH40 mem_exe_result_reg_29_ ( .D(n172), .CK(clk), .Q(
        mem_exe_result[29]) );
  DQV4_8TH40 mem_exe_result_reg_28_ ( .D(n171), .CK(clk), .Q(
        mem_exe_result[28]) );
  DQV4_8TH40 mem_exe_result_reg_27_ ( .D(n170), .CK(clk), .Q(
        mem_exe_result[27]) );
  DQV4_8TH40 mem_exe_result_reg_26_ ( .D(n169), .CK(clk), .Q(
        mem_exe_result[26]) );
  DQV4_8TH40 mem_exe_result_reg_25_ ( .D(n168), .CK(clk), .Q(
        mem_exe_result[25]) );
  DQV4_8TH40 mem_exe_result_reg_24_ ( .D(n167), .CK(clk), .Q(
        mem_exe_result[24]) );
  DQV4_8TH40 mem_exe_result_reg_23_ ( .D(n166), .CK(clk), .Q(
        mem_exe_result[23]) );
  DQV4_8TH40 mem_exe_result_reg_22_ ( .D(n165), .CK(clk), .Q(
        mem_exe_result[22]) );
  DQV4_8TH40 mem_exe_result_reg_21_ ( .D(n164), .CK(clk), .Q(
        mem_exe_result[21]) );
  DQV4_8TH40 mem_exe_result_reg_20_ ( .D(n163), .CK(clk), .Q(
        mem_exe_result[20]) );
  DQV4_8TH40 mem_exe_result_reg_19_ ( .D(n162), .CK(clk), .Q(
        mem_exe_result[19]) );
  DQV4_8TH40 mem_exe_result_reg_18_ ( .D(n161), .CK(clk), .Q(
        mem_exe_result[18]) );
  DQV4_8TH40 mem_exe_result_reg_17_ ( .D(n160), .CK(clk), .Q(
        mem_exe_result[17]) );
  DQV4_8TH40 mem_exe_result_reg_16_ ( .D(n159), .CK(clk), .Q(
        mem_exe_result[16]) );
  DQV4_8TH40 mem_exe_result_reg_15_ ( .D(n158), .CK(clk), .Q(
        mem_exe_result[15]) );
  DQV4_8TH40 mem_exe_result_reg_14_ ( .D(n157), .CK(clk), .Q(
        mem_exe_result[14]) );
  DQV4_8TH40 mem_exe_result_reg_13_ ( .D(n156), .CK(clk), .Q(
        mem_exe_result[13]) );
  DQV4_8TH40 mem_exe_result_reg_12_ ( .D(n155), .CK(clk), .Q(
        mem_exe_result[12]) );
  DQV4_8TH40 mem_exe_result_reg_11_ ( .D(n154), .CK(clk), .Q(
        mem_exe_result[11]) );
  DQV4_8TH40 mem_exe_result_reg_10_ ( .D(n153), .CK(clk), .Q(
        mem_exe_result[10]) );
  DQV4_8TH40 mem_exe_result_reg_9_ ( .D(n152), .CK(clk), .Q(mem_exe_result[9])
         );
  DQV4_8TH40 mem_exe_result_reg_8_ ( .D(n151), .CK(clk), .Q(mem_exe_result[8])
         );
  DQV4_8TH40 mem_exe_result_reg_7_ ( .D(n150), .CK(clk), .Q(mem_exe_result[7])
         );
  DQV4_8TH40 mem_exe_result_reg_6_ ( .D(n149), .CK(clk), .Q(mem_exe_result[6])
         );
  DQV4_8TH40 mem_exe_result_reg_5_ ( .D(n148), .CK(clk), .Q(mem_exe_result[5])
         );
  DQV4_8TH40 mem_exe_result_reg_4_ ( .D(n147), .CK(clk), .Q(mem_exe_result[4])
         );
  DQV4_8TH40 mem_exe_result_reg_3_ ( .D(n146), .CK(clk), .Q(mem_exe_result[3])
         );
  DQV4_8TH40 mem_exe_result_reg_2_ ( .D(n145), .CK(clk), .Q(mem_exe_result[2])
         );
  DQV4_8TH40 mem_exe_result_reg_1_ ( .D(n144), .CK(clk), .Q(mem_exe_result[1])
         );
  DQV4_8TH40 mem_exe_result_reg_0_ ( .D(n143), .CK(clk), .Q(mem_exe_result[0])
         );
  DQV4_8TH40 mem_hi_reg_31_ ( .D(n142), .CK(clk), .Q(mem_hi[31]) );
  DQV4_8TH40 mem_hi_reg_30_ ( .D(n141), .CK(clk), .Q(mem_hi[30]) );
  DQV4_8TH40 mem_hi_reg_29_ ( .D(n140), .CK(clk), .Q(mem_hi[29]) );
  DQV4_8TH40 mem_hi_reg_28_ ( .D(n139), .CK(clk), .Q(mem_hi[28]) );
  DQV4_8TH40 mem_hi_reg_27_ ( .D(n138), .CK(clk), .Q(mem_hi[27]) );
  DQV4_8TH40 mem_hi_reg_26_ ( .D(n137), .CK(clk), .Q(mem_hi[26]) );
  DQV4_8TH40 mem_hi_reg_25_ ( .D(n136), .CK(clk), .Q(mem_hi[25]) );
  DQV4_8TH40 mem_hi_reg_24_ ( .D(n135), .CK(clk), .Q(mem_hi[24]) );
  DQV4_8TH40 mem_hi_reg_23_ ( .D(n134), .CK(clk), .Q(mem_hi[23]) );
  DQV4_8TH40 mem_hi_reg_22_ ( .D(n133), .CK(clk), .Q(mem_hi[22]) );
  DQV4_8TH40 mem_hi_reg_21_ ( .D(n132), .CK(clk), .Q(mem_hi[21]) );
  DQV4_8TH40 mem_hi_reg_20_ ( .D(n131), .CK(clk), .Q(mem_hi[20]) );
  DQV4_8TH40 mem_hi_reg_19_ ( .D(n130), .CK(clk), .Q(mem_hi[19]) );
  DQV4_8TH40 mem_hi_reg_18_ ( .D(n129), .CK(clk), .Q(mem_hi[18]) );
  DQV4_8TH40 mem_hi_reg_17_ ( .D(n128), .CK(clk), .Q(mem_hi[17]) );
  DQV4_8TH40 mem_hi_reg_16_ ( .D(n127), .CK(clk), .Q(mem_hi[16]) );
  DQV4_8TH40 mem_hi_reg_15_ ( .D(n126), .CK(clk), .Q(mem_hi[15]) );
  DQV4_8TH40 mem_hi_reg_14_ ( .D(n125), .CK(clk), .Q(mem_hi[14]) );
  DQV4_8TH40 mem_hi_reg_13_ ( .D(n124), .CK(clk), .Q(mem_hi[13]) );
  DQV4_8TH40 mem_hi_reg_12_ ( .D(n123), .CK(clk), .Q(mem_hi[12]) );
  DQV4_8TH40 mem_hi_reg_11_ ( .D(n122), .CK(clk), .Q(mem_hi[11]) );
  DQV4_8TH40 mem_hi_reg_10_ ( .D(n121), .CK(clk), .Q(mem_hi[10]) );
  DQV4_8TH40 mem_hi_reg_9_ ( .D(n120), .CK(clk), .Q(mem_hi[9]) );
  DQV4_8TH40 mem_hi_reg_8_ ( .D(n119), .CK(clk), .Q(mem_hi[8]) );
  DQV4_8TH40 mem_hi_reg_7_ ( .D(n118), .CK(clk), .Q(mem_hi[7]) );
  DQV4_8TH40 mem_hi_reg_6_ ( .D(n117), .CK(clk), .Q(mem_hi[6]) );
  DQV4_8TH40 mem_hi_reg_5_ ( .D(n116), .CK(clk), .Q(mem_hi[5]) );
  DQV4_8TH40 mem_hi_reg_4_ ( .D(n115), .CK(clk), .Q(mem_hi[4]) );
  DQV4_8TH40 mem_hi_reg_3_ ( .D(n114), .CK(clk), .Q(mem_hi[3]) );
  DQV4_8TH40 mem_hi_reg_2_ ( .D(n113), .CK(clk), .Q(mem_hi[2]) );
  DQV4_8TH40 mem_hi_reg_1_ ( .D(n112), .CK(clk), .Q(mem_hi[1]) );
  DQV4_8TH40 mem_hi_reg_0_ ( .D(n111), .CK(clk), .Q(mem_hi[0]) );
  DQV4_8TH40 mem_lo_reg_31_ ( .D(n110), .CK(clk), .Q(mem_lo[31]) );
  DQV4_8TH40 mem_lo_reg_30_ ( .D(n109), .CK(clk), .Q(mem_lo[30]) );
  DQV4_8TH40 mem_lo_reg_29_ ( .D(n108), .CK(clk), .Q(mem_lo[29]) );
  DQV4_8TH40 mem_lo_reg_28_ ( .D(n107), .CK(clk), .Q(mem_lo[28]) );
  DQV4_8TH40 mem_lo_reg_27_ ( .D(n106), .CK(clk), .Q(mem_lo[27]) );
  DQV4_8TH40 mem_lo_reg_26_ ( .D(n105), .CK(clk), .Q(mem_lo[26]) );
  DQV4_8TH40 mem_lo_reg_25_ ( .D(n104), .CK(clk), .Q(mem_lo[25]) );
  DQV4_8TH40 mem_lo_reg_24_ ( .D(n103), .CK(clk), .Q(mem_lo[24]) );
  DQV4_8TH40 mem_lo_reg_23_ ( .D(n102), .CK(clk), .Q(mem_lo[23]) );
  DQV4_8TH40 mem_lo_reg_22_ ( .D(n101), .CK(clk), .Q(mem_lo[22]) );
  DQV4_8TH40 mem_lo_reg_21_ ( .D(n100), .CK(clk), .Q(mem_lo[21]) );
  DQV4_8TH40 mem_lo_reg_20_ ( .D(n99), .CK(clk), .Q(mem_lo[20]) );
  DQV4_8TH40 mem_lo_reg_19_ ( .D(n98), .CK(clk), .Q(mem_lo[19]) );
  DQV4_8TH40 mem_lo_reg_18_ ( .D(n97), .CK(clk), .Q(mem_lo[18]) );
  DQV4_8TH40 mem_lo_reg_17_ ( .D(n96), .CK(clk), .Q(mem_lo[17]) );
  DQV4_8TH40 mem_lo_reg_16_ ( .D(n95), .CK(clk), .Q(mem_lo[16]) );
  DQV4_8TH40 mem_lo_reg_15_ ( .D(n94), .CK(clk), .Q(mem_lo[15]) );
  DQV4_8TH40 mem_lo_reg_14_ ( .D(n93), .CK(clk), .Q(mem_lo[14]) );
  DQV4_8TH40 mem_lo_reg_13_ ( .D(n92), .CK(clk), .Q(mem_lo[13]) );
  DQV4_8TH40 mem_lo_reg_12_ ( .D(n91), .CK(clk), .Q(mem_lo[12]) );
  DQV4_8TH40 mem_lo_reg_11_ ( .D(n90), .CK(clk), .Q(mem_lo[11]) );
  DQV4_8TH40 mem_lo_reg_10_ ( .D(n89), .CK(clk), .Q(mem_lo[10]) );
  DQV4_8TH40 mem_lo_reg_9_ ( .D(n88), .CK(clk), .Q(mem_lo[9]) );
  DQV4_8TH40 mem_lo_reg_8_ ( .D(n87), .CK(clk), .Q(mem_lo[8]) );
  DQV4_8TH40 mem_lo_reg_7_ ( .D(n86), .CK(clk), .Q(mem_lo[7]) );
  DQV4_8TH40 mem_lo_reg_6_ ( .D(n85), .CK(clk), .Q(mem_lo[6]) );
  DQV4_8TH40 mem_lo_reg_5_ ( .D(n84), .CK(clk), .Q(mem_lo[5]) );
  DQV4_8TH40 mem_lo_reg_4_ ( .D(n83), .CK(clk), .Q(mem_lo[4]) );
  DQV4_8TH40 mem_lo_reg_3_ ( .D(n82), .CK(clk), .Q(mem_lo[3]) );
  DQV4_8TH40 mem_lo_reg_2_ ( .D(n81), .CK(clk), .Q(mem_lo[2]) );
  DQV4_8TH40 mem_lo_reg_1_ ( .D(n80), .CK(clk), .Q(mem_lo[1]) );
  DQV4_8TH40 mem_lo_reg_0_ ( .D(n79), .CK(clk), .Q(mem_lo[0]) );
  DQV4_8TH40 mem_hilo_we_reg ( .D(n78), .CK(clk), .Q(mem_hilo_we) );
  DQV4_8TH40 mem_inst_type_reg_7_ ( .D(n77), .CK(clk), .Q(mem_inst_type[7]) );
  DQV4_8TH40 mem_inst_type_reg_6_ ( .D(n76), .CK(clk), .Q(mem_inst_type[6]) );
  DQV4_8TH40 mem_inst_type_reg_5_ ( .D(n75), .CK(clk), .Q(mem_inst_type[5]) );
  DQV4_8TH40 mem_inst_type_reg_4_ ( .D(n74), .CK(clk), .Q(mem_inst_type[4]) );
  DQV4_8TH40 mem_inst_type_reg_3_ ( .D(n73), .CK(clk), .Q(mem_inst_type[3]) );
  DQV4_8TH40 mem_inst_type_reg_2_ ( .D(n72), .CK(clk), .Q(mem_inst_type[2]) );
  DQV4_8TH40 mem_inst_type_reg_1_ ( .D(n71), .CK(clk), .Q(mem_inst_type[1]) );
  DQV4_8TH40 mem_inst_type_reg_0_ ( .D(n70), .CK(clk), .Q(mem_inst_type[0]) );
  DQV4_8TH40 mem_dmem_addr_reg_31_ ( .D(n69), .CK(clk), .Q(mem_dmem_addr[31])
         );
  DQV4_8TH40 mem_dmem_addr_reg_30_ ( .D(n68), .CK(clk), .Q(mem_dmem_addr[30])
         );
  DQV4_8TH40 mem_dmem_addr_reg_29_ ( .D(n67), .CK(clk), .Q(mem_dmem_addr[29])
         );
  DQV4_8TH40 mem_dmem_addr_reg_28_ ( .D(n66), .CK(clk), .Q(mem_dmem_addr[28])
         );
  DQV4_8TH40 mem_dmem_addr_reg_27_ ( .D(n65), .CK(clk), .Q(mem_dmem_addr[27])
         );
  DQV4_8TH40 mem_dmem_addr_reg_26_ ( .D(n64), .CK(clk), .Q(mem_dmem_addr[26])
         );
  DQV4_8TH40 mem_dmem_addr_reg_25_ ( .D(n63), .CK(clk), .Q(mem_dmem_addr[25])
         );
  DQV4_8TH40 mem_dmem_addr_reg_24_ ( .D(n62), .CK(clk), .Q(mem_dmem_addr[24])
         );
  DQV4_8TH40 mem_dmem_addr_reg_23_ ( .D(n61), .CK(clk), .Q(mem_dmem_addr[23])
         );
  DQV4_8TH40 mem_dmem_addr_reg_22_ ( .D(n60), .CK(clk), .Q(mem_dmem_addr[22])
         );
  DQV4_8TH40 mem_dmem_addr_reg_21_ ( .D(n59), .CK(clk), .Q(mem_dmem_addr[21])
         );
  DQV4_8TH40 mem_dmem_addr_reg_20_ ( .D(n58), .CK(clk), .Q(mem_dmem_addr[20])
         );
  DQV4_8TH40 mem_dmem_addr_reg_19_ ( .D(n57), .CK(clk), .Q(mem_dmem_addr[19])
         );
  DQV4_8TH40 mem_dmem_addr_reg_18_ ( .D(n56), .CK(clk), .Q(mem_dmem_addr[18])
         );
  DQV4_8TH40 mem_dmem_addr_reg_17_ ( .D(n55), .CK(clk), .Q(mem_dmem_addr[17])
         );
  DQV4_8TH40 mem_dmem_addr_reg_16_ ( .D(n54), .CK(clk), .Q(mem_dmem_addr[16])
         );
  DQV4_8TH40 mem_dmem_addr_reg_15_ ( .D(n53), .CK(clk), .Q(mem_dmem_addr[15])
         );
  DQV4_8TH40 mem_dmem_addr_reg_14_ ( .D(n52), .CK(clk), .Q(mem_dmem_addr[14])
         );
  DQV4_8TH40 mem_dmem_addr_reg_13_ ( .D(n51), .CK(clk), .Q(mem_dmem_addr[13])
         );
  DQV4_8TH40 mem_dmem_addr_reg_12_ ( .D(n50), .CK(clk), .Q(mem_dmem_addr[12])
         );
  DQV4_8TH40 mem_dmem_addr_reg_11_ ( .D(n49), .CK(clk), .Q(mem_dmem_addr[11])
         );
  DQV4_8TH40 mem_dmem_addr_reg_10_ ( .D(n48), .CK(clk), .Q(mem_dmem_addr[10])
         );
  DQV4_8TH40 mem_dmem_addr_reg_9_ ( .D(n47), .CK(clk), .Q(mem_dmem_addr[9]) );
  DQV4_8TH40 mem_dmem_addr_reg_8_ ( .D(n46), .CK(clk), .Q(mem_dmem_addr[8]) );
  DQV4_8TH40 mem_dmem_addr_reg_7_ ( .D(n45), .CK(clk), .Q(mem_dmem_addr[7]) );
  DQV4_8TH40 mem_dmem_addr_reg_6_ ( .D(n44), .CK(clk), .Q(mem_dmem_addr[6]) );
  DQV4_8TH40 mem_dmem_addr_reg_5_ ( .D(n43), .CK(clk), .Q(mem_dmem_addr[5]) );
  DQV4_8TH40 mem_dmem_addr_reg_4_ ( .D(n42), .CK(clk), .Q(mem_dmem_addr[4]) );
  DQV4_8TH40 mem_dmem_addr_reg_3_ ( .D(n41), .CK(clk), .Q(mem_dmem_addr[3]) );
  DQV4_8TH40 mem_dmem_addr_reg_2_ ( .D(n40), .CK(clk), .Q(mem_dmem_addr[2]) );
  DQV4_8TH40 mem_dmem_addr_reg_1_ ( .D(n39), .CK(clk), .Q(mem_dmem_addr[1]) );
  DQV4_8TH40 mem_dmem_addr_reg_0_ ( .D(n38), .CK(clk), .Q(mem_dmem_addr[0]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_31_ ( .D(n37), .CK(clk), .Q(
        mem_ls_data_tmp[31]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_30_ ( .D(n36), .CK(clk), .Q(
        mem_ls_data_tmp[30]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_29_ ( .D(n35), .CK(clk), .Q(
        mem_ls_data_tmp[29]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_28_ ( .D(n34), .CK(clk), .Q(
        mem_ls_data_tmp[28]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_27_ ( .D(n33), .CK(clk), .Q(
        mem_ls_data_tmp[27]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_26_ ( .D(n32), .CK(clk), .Q(
        mem_ls_data_tmp[26]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_25_ ( .D(n31), .CK(clk), .Q(
        mem_ls_data_tmp[25]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_24_ ( .D(n30), .CK(clk), .Q(
        mem_ls_data_tmp[24]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_23_ ( .D(n29), .CK(clk), .Q(
        mem_ls_data_tmp[23]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_22_ ( .D(n28), .CK(clk), .Q(
        mem_ls_data_tmp[22]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_21_ ( .D(n27), .CK(clk), .Q(
        mem_ls_data_tmp[21]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_20_ ( .D(n26), .CK(clk), .Q(
        mem_ls_data_tmp[20]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_19_ ( .D(n25), .CK(clk), .Q(
        mem_ls_data_tmp[19]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_18_ ( .D(n24), .CK(clk), .Q(
        mem_ls_data_tmp[18]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_17_ ( .D(n23), .CK(clk), .Q(
        mem_ls_data_tmp[17]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_16_ ( .D(n22), .CK(clk), .Q(
        mem_ls_data_tmp[16]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_15_ ( .D(n21), .CK(clk), .Q(
        mem_ls_data_tmp[15]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_14_ ( .D(n20), .CK(clk), .Q(
        mem_ls_data_tmp[14]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_13_ ( .D(n19), .CK(clk), .Q(
        mem_ls_data_tmp[13]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_12_ ( .D(n18), .CK(clk), .Q(
        mem_ls_data_tmp[12]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_11_ ( .D(n17), .CK(clk), .Q(
        mem_ls_data_tmp[11]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_10_ ( .D(n16), .CK(clk), .Q(
        mem_ls_data_tmp[10]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_9_ ( .D(n15), .CK(clk), .Q(mem_ls_data_tmp[9]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_8_ ( .D(n14), .CK(clk), .Q(mem_ls_data_tmp[8]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_7_ ( .D(n13), .CK(clk), .Q(mem_ls_data_tmp[7]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_6_ ( .D(n12), .CK(clk), .Q(mem_ls_data_tmp[6]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_5_ ( .D(n11), .CK(clk), .Q(mem_ls_data_tmp[5]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_4_ ( .D(n10), .CK(clk), .Q(mem_ls_data_tmp[4]) );
  DQV4_8TH40 mem_ls_data_tmp_reg_3_ ( .D(n9), .CK(clk), .Q(mem_ls_data_tmp[3])
         );
  DQV4_8TH40 mem_ls_data_tmp_reg_2_ ( .D(n8), .CK(clk), .Q(mem_ls_data_tmp[2])
         );
  DQV4_8TH40 mem_ls_data_tmp_reg_1_ ( .D(n7), .CK(clk), .Q(mem_ls_data_tmp[1])
         );
  DQV4_8TH40 mem_ls_data_tmp_reg_0_ ( .D(n6), .CK(clk), .Q(mem_ls_data_tmp[0])
         );
  DQV4_8TH40 mem_cp0_we_reg ( .D(n5), .CK(clk), .Q(mem_cp0_we) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_63_ ( .D(ex_hilo_tmp_i[63]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[63]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_62_ ( .D(ex_hilo_tmp_i[62]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[62]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_61_ ( .D(ex_hilo_tmp_i[61]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[61]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_60_ ( .D(ex_hilo_tmp_i[60]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[60]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_59_ ( .D(ex_hilo_tmp_i[59]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[59]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_58_ ( .D(ex_hilo_tmp_i[58]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[58]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_57_ ( .D(ex_hilo_tmp_i[57]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[57]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_56_ ( .D(ex_hilo_tmp_i[56]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[56]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_55_ ( .D(ex_hilo_tmp_i[55]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[55]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_54_ ( .D(ex_hilo_tmp_i[54]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[54]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_53_ ( .D(ex_hilo_tmp_i[53]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[53]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_52_ ( .D(ex_hilo_tmp_i[52]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[52]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_51_ ( .D(ex_hilo_tmp_i[51]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[51]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_50_ ( .D(ex_hilo_tmp_i[50]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[50]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_49_ ( .D(ex_hilo_tmp_i[49]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[49]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_48_ ( .D(ex_hilo_tmp_i[48]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[48]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_47_ ( .D(ex_hilo_tmp_i[47]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[47]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_46_ ( .D(ex_hilo_tmp_i[46]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[46]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_45_ ( .D(ex_hilo_tmp_i[45]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[45]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_44_ ( .D(ex_hilo_tmp_i[44]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[44]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_43_ ( .D(ex_hilo_tmp_i[43]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[43]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_42_ ( .D(ex_hilo_tmp_i[42]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[42]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_41_ ( .D(ex_hilo_tmp_i[41]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[41]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_40_ ( .D(ex_hilo_tmp_i[40]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[40]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_39_ ( .D(ex_hilo_tmp_i[39]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[39]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_38_ ( .D(ex_hilo_tmp_i[38]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[38]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_37_ ( .D(ex_hilo_tmp_i[37]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[37]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_36_ ( .D(ex_hilo_tmp_i[36]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[36]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_35_ ( .D(ex_hilo_tmp_i[35]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[35]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_34_ ( .D(ex_hilo_tmp_i[34]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[34]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_33_ ( .D(ex_hilo_tmp_i[33]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[33]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_32_ ( .D(ex_hilo_tmp_i[32]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[32]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_31_ ( .D(ex_hilo_tmp_i[31]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[31]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_30_ ( .D(ex_hilo_tmp_i[30]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[30]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_29_ ( .D(ex_hilo_tmp_i[29]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[29]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_28_ ( .D(ex_hilo_tmp_i[28]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[28]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_27_ ( .D(ex_hilo_tmp_i[27]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[27]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_26_ ( .D(ex_hilo_tmp_i[26]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[26]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_25_ ( .D(ex_hilo_tmp_i[25]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[25]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_24_ ( .D(ex_hilo_tmp_i[24]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[24]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_23_ ( .D(ex_hilo_tmp_i[23]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[23]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_22_ ( .D(ex_hilo_tmp_i[22]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[22]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_21_ ( .D(ex_hilo_tmp_i[21]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[21]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_20_ ( .D(ex_hilo_tmp_i[20]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[20]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_19_ ( .D(ex_hilo_tmp_i[19]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[19]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_18_ ( .D(ex_hilo_tmp_i[18]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[18]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_17_ ( .D(ex_hilo_tmp_i[17]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[17]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_16_ ( .D(ex_hilo_tmp_i[16]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[16]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_15_ ( .D(ex_hilo_tmp_i[15]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[15]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_14_ ( .D(ex_hilo_tmp_i[14]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[14]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_13_ ( .D(ex_hilo_tmp_i[13]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[13]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_12_ ( .D(ex_hilo_tmp_i[12]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[12]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_11_ ( .D(ex_hilo_tmp_i[11]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[11]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_10_ ( .D(ex_hilo_tmp_i[10]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[10]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_9_ ( .D(ex_hilo_tmp_i[9]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[9]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_8_ ( .D(ex_hilo_tmp_i[8]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[8]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_7_ ( .D(ex_hilo_tmp_i[7]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[7]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_6_ ( .D(ex_hilo_tmp_i[6]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[6]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_5_ ( .D(ex_hilo_tmp_i[5]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[5]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_4_ ( .D(ex_hilo_tmp_i[4]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[4]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_3_ ( .D(ex_hilo_tmp_i[3]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[3]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_2_ ( .D(ex_hilo_tmp_i[2]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[2]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_1_ ( .D(ex_hilo_tmp_i[1]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[1]) );
  DGRNQV4_8TH40 ex_hilo_tmp_o_reg_0_ ( .D(ex_hilo_tmp_i[0]), .RN(n313), .CK(
        clk), .Q(ex_hilo_tmp_o[0]) );
  DGRNQV4_8TH40 ex_cycl_cnt_o_reg_1_ ( .D(ex_cycl_cnt_i[1]), .RN(n313), .CK(
        clk), .Q(ex_cycl_cnt_o[1]) );
  DGRNQV4_8TH40 ex_cycl_cnt_o_reg_0_ ( .D(ex_cycl_cnt_i[0]), .RN(n313), .CK(
        clk), .Q(ex_cycl_cnt_o[0]) );
  NAND2V2_8TH40 U3 ( .A1(stall_ctrl[4]), .A2(n313), .ZN(n1) );
  AO22V4_8TH40 U4 ( .A1(mem_hilo_we), .A2(n226), .B1(ex_hilo_we), .B2(n288), 
        .Z(n78) );
  AO22V4_8TH40 U5 ( .A1(mem_lo[0]), .A2(n222), .B1(ex_lo[0]), .B2(n289), .Z(
        n79) );
  AO22V4_8TH40 U6 ( .A1(mem_lo[1]), .A2(n219), .B1(ex_lo[1]), .B2(n289), .Z(
        n80) );
  AO22V4_8TH40 U7 ( .A1(mem_lo[2]), .A2(n220), .B1(ex_lo[2]), .B2(n289), .Z(
        n81) );
  AO22V4_8TH40 U8 ( .A1(mem_lo[3]), .A2(n221), .B1(ex_lo[3]), .B2(n289), .Z(
        n82) );
  AO22V4_8TH40 U9 ( .A1(mem_lo[4]), .A2(n232), .B1(ex_lo[4]), .B2(n289), .Z(
        n83) );
  AO22V4_8TH40 U10 ( .A1(mem_lo[5]), .A2(n236), .B1(ex_lo[5]), .B2(n289), .Z(
        n84) );
  AO22V4_8TH40 U11 ( .A1(mem_lo[6]), .A2(n236), .B1(ex_lo[6]), .B2(n289), .Z(
        n85) );
  AO22V4_8TH40 U12 ( .A1(mem_lo[7]), .A2(n236), .B1(ex_lo[7]), .B2(n289), .Z(
        n86) );
  AO22V4_8TH40 U13 ( .A1(mem_lo[8]), .A2(n236), .B1(ex_lo[8]), .B2(n289), .Z(
        n87) );
  AO22V4_8TH40 U14 ( .A1(mem_lo[9]), .A2(n236), .B1(ex_lo[9]), .B2(n289), .Z(
        n88) );
  AO22V4_8TH40 U15 ( .A1(mem_lo[10]), .A2(n236), .B1(ex_lo[10]), .B2(n289), 
        .Z(n89) );
  AO22V4_8TH40 U16 ( .A1(mem_lo[11]), .A2(n236), .B1(ex_lo[11]), .B2(n290), 
        .Z(n90) );
  AO22V4_8TH40 U17 ( .A1(mem_lo[12]), .A2(n236), .B1(ex_lo[12]), .B2(n290), 
        .Z(n91) );
  AO22V4_8TH40 U18 ( .A1(mem_lo[13]), .A2(n236), .B1(ex_lo[13]), .B2(n290), 
        .Z(n92) );
  AO22V4_8TH40 U19 ( .A1(mem_lo[14]), .A2(n236), .B1(ex_lo[14]), .B2(n290), 
        .Z(n93) );
  AO22V4_8TH40 U20 ( .A1(mem_lo[15]), .A2(n236), .B1(ex_lo[15]), .B2(n290), 
        .Z(n94) );
  AO22V4_8TH40 U21 ( .A1(mem_lo[16]), .A2(n236), .B1(ex_lo[16]), .B2(n290), 
        .Z(n95) );
  AO22V4_8TH40 U22 ( .A1(mem_lo[17]), .A2(n232), .B1(ex_lo[17]), .B2(n290), 
        .Z(n96) );
  AO22V4_8TH40 U23 ( .A1(mem_lo[18]), .A2(n233), .B1(ex_lo[18]), .B2(n290), 
        .Z(n97) );
  AO22V4_8TH40 U24 ( .A1(mem_lo[19]), .A2(n220), .B1(ex_lo[19]), .B2(n290), 
        .Z(n98) );
  AO22V4_8TH40 U25 ( .A1(mem_lo[20]), .A2(n221), .B1(ex_lo[20]), .B2(n290), 
        .Z(n99) );
  AO22V4_8TH40 U26 ( .A1(mem_lo[21]), .A2(n2), .B1(ex_lo[21]), .B2(n247), .Z(
        n100) );
  AO22V4_8TH40 U27 ( .A1(mem_lo[22]), .A2(n2), .B1(ex_lo[22]), .B2(n247), .Z(
        n101) );
  AO22V4_8TH40 U28 ( .A1(mem_lo[23]), .A2(n2), .B1(ex_lo[23]), .B2(n247), .Z(
        n102) );
  AO22V4_8TH40 U29 ( .A1(mem_lo[24]), .A2(n2), .B1(ex_lo[24]), .B2(n247), .Z(
        n103) );
  AO22V4_8TH40 U30 ( .A1(mem_lo[25]), .A2(n2), .B1(ex_lo[25]), .B2(n247), .Z(
        n104) );
  AO22V4_8TH40 U31 ( .A1(mem_lo[26]), .A2(n2), .B1(ex_lo[26]), .B2(n247), .Z(
        n105) );
  AO22V4_8TH40 U32 ( .A1(mem_lo[27]), .A2(n2), .B1(ex_lo[27]), .B2(n247), .Z(
        n106) );
  AO22V4_8TH40 U33 ( .A1(mem_lo[28]), .A2(n2), .B1(ex_lo[28]), .B2(n247), .Z(
        n107) );
  AO22V4_8TH40 U34 ( .A1(mem_lo[29]), .A2(n2), .B1(ex_lo[29]), .B2(n247), .Z(
        n108) );
  AO22V4_8TH40 U35 ( .A1(mem_lo[30]), .A2(n2), .B1(ex_lo[30]), .B2(n247), .Z(
        n109) );
  AO22V4_8TH40 U36 ( .A1(mem_lo[31]), .A2(n2), .B1(ex_lo[31]), .B2(n248), .Z(
        n110) );
  AO22V4_8TH40 U37 ( .A1(mem_hi[0]), .A2(n3), .B1(ex_hi[0]), .B2(n248), .Z(
        n111) );
  AO22V4_8TH40 U38 ( .A1(mem_hi[1]), .A2(n3), .B1(ex_hi[1]), .B2(n248), .Z(
        n112) );
  AO22V4_8TH40 U39 ( .A1(mem_hi[2]), .A2(n3), .B1(ex_hi[2]), .B2(n248), .Z(
        n113) );
  AO22V4_8TH40 U40 ( .A1(mem_hi[3]), .A2(n3), .B1(ex_hi[3]), .B2(n248), .Z(
        n114) );
  AO22V4_8TH40 U41 ( .A1(mem_hi[4]), .A2(n3), .B1(ex_hi[4]), .B2(n248), .Z(
        n115) );
  AO22V4_8TH40 U42 ( .A1(mem_hi[5]), .A2(n3), .B1(ex_hi[5]), .B2(n248), .Z(
        n116) );
  AO22V4_8TH40 U43 ( .A1(mem_hi[6]), .A2(n3), .B1(ex_hi[6]), .B2(n248), .Z(
        n117) );
  AO22V4_8TH40 U44 ( .A1(mem_hi[7]), .A2(n3), .B1(ex_hi[7]), .B2(n248), .Z(
        n118) );
  AO22V4_8TH40 U45 ( .A1(mem_hi[8]), .A2(n3), .B1(ex_hi[8]), .B2(n248), .Z(
        n119) );
  AO22V4_8TH40 U46 ( .A1(mem_hi[9]), .A2(n3), .B1(ex_hi[9]), .B2(n248), .Z(
        n120) );
  AO22V4_8TH40 U47 ( .A1(mem_hi[10]), .A2(n3), .B1(ex_hi[10]), .B2(n283), .Z(
        n121) );
  AO22V4_8TH40 U48 ( .A1(mem_hi[11]), .A2(n3), .B1(ex_hi[11]), .B2(n249), .Z(
        n122) );
  AO22V4_8TH40 U49 ( .A1(mem_hi[12]), .A2(n4), .B1(ex_hi[12]), .B2(n285), .Z(
        n123) );
  AO22V4_8TH40 U50 ( .A1(mem_hi[13]), .A2(n4), .B1(ex_hi[13]), .B2(n288), .Z(
        n124) );
  AO22V4_8TH40 U51 ( .A1(mem_hi[14]), .A2(n4), .B1(ex_hi[14]), .B2(n312), .Z(
        n125) );
  AO22V4_8TH40 U52 ( .A1(mem_hi[15]), .A2(n4), .B1(ex_hi[15]), .B2(n290), .Z(
        n126) );
  AO22V4_8TH40 U53 ( .A1(mem_hi[16]), .A2(n4), .B1(ex_hi[16]), .B2(n283), .Z(
        n127) );
  AO22V4_8TH40 U54 ( .A1(mem_hi[17]), .A2(n4), .B1(ex_hi[17]), .B2(n284), .Z(
        n128) );
  AO22V4_8TH40 U55 ( .A1(mem_hi[18]), .A2(n4), .B1(ex_hi[18]), .B2(n247), .Z(
        n129) );
  AO22V4_8TH40 U56 ( .A1(mem_hi[19]), .A2(n4), .B1(ex_hi[19]), .B2(n248), .Z(
        n130) );
  AO22V4_8TH40 U57 ( .A1(mem_hi[20]), .A2(n4), .B1(ex_hi[20]), .B2(n286), .Z(
        n131) );
  AO22V4_8TH40 U58 ( .A1(mem_hi[21]), .A2(n4), .B1(ex_hi[21]), .B2(n249), .Z(
        n132) );
  AO22V4_8TH40 U59 ( .A1(mem_hi[22]), .A2(n4), .B1(ex_hi[22]), .B2(n249), .Z(
        n133) );
  AO22V4_8TH40 U60 ( .A1(mem_hi[23]), .A2(n4), .B1(ex_hi[23]), .B2(n249), .Z(
        n134) );
  AO22V4_8TH40 U61 ( .A1(mem_hi[24]), .A2(n219), .B1(ex_hi[24]), .B2(n249), 
        .Z(n135) );
  AO22V4_8TH40 U62 ( .A1(mem_hi[25]), .A2(n219), .B1(ex_hi[25]), .B2(n249), 
        .Z(n136) );
  AO22V4_8TH40 U63 ( .A1(mem_hi[26]), .A2(n219), .B1(ex_hi[26]), .B2(n249), 
        .Z(n137) );
  AO22V4_8TH40 U64 ( .A1(mem_hi[27]), .A2(n219), .B1(ex_hi[27]), .B2(n249), 
        .Z(n138) );
  AO22V4_8TH40 U65 ( .A1(mem_hi[28]), .A2(n219), .B1(ex_hi[28]), .B2(n249), 
        .Z(n139) );
  AO22V4_8TH40 U66 ( .A1(mem_hi[29]), .A2(n219), .B1(ex_hi[29]), .B2(n249), 
        .Z(n140) );
  AO22V4_8TH40 U67 ( .A1(mem_hi[30]), .A2(n219), .B1(ex_hi[30]), .B2(n249), 
        .Z(n141) );
  AO22V4_8TH40 U68 ( .A1(mem_hi[31]), .A2(n219), .B1(ex_hi[31]), .B2(n249), 
        .Z(n142) );
  AO22V4_8TH40 U69 ( .A1(mem_cp0_waddr[0]), .A2(n225), .B1(ex_cp0_waddr[0]), 
        .B2(n284), .Z(n214) );
  AO22V4_8TH40 U70 ( .A1(mem_cp0_waddr[1]), .A2(n225), .B1(ex_cp0_waddr[1]), 
        .B2(n284), .Z(n215) );
  AO22V4_8TH40 U71 ( .A1(mem_except_type[10]), .A2(n226), .B1(
        ex_except_type[10]), .B2(n250), .Z(n229) );
  AO22V4_8TH40 U72 ( .A1(mem_cp0_wdata[0]), .A2(n223), .B1(ex_cp0_wdata[0]), 
        .B2(n250), .Z(n182) );
  AO22V4_8TH40 U73 ( .A1(mem_cp0_wdata[1]), .A2(n223), .B1(ex_cp0_wdata[1]), 
        .B2(n285), .Z(n183) );
  AO22V4_8TH40 U74 ( .A1(mem_cp0_wdata[2]), .A2(n223), .B1(ex_cp0_wdata[2]), 
        .B2(n286), .Z(n184) );
  AO22V4_8TH40 U75 ( .A1(mem_cp0_wdata[3]), .A2(n223), .B1(ex_cp0_wdata[3]), 
        .B2(n286), .Z(n185) );
  AO22V4_8TH40 U76 ( .A1(mem_cp0_wdata[4]), .A2(n223), .B1(ex_cp0_wdata[4]), 
        .B2(n288), .Z(n186) );
  AO22V4_8TH40 U77 ( .A1(mem_cp0_wdata[5]), .A2(n223), .B1(ex_cp0_wdata[5]), 
        .B2(n283), .Z(n187) );
  AO22V4_8TH40 U78 ( .A1(mem_cp0_wdata[6]), .A2(n223), .B1(ex_cp0_wdata[6]), 
        .B2(n283), .Z(n188) );
  AO22V4_8TH40 U79 ( .A1(mem_cp0_wdata[7]), .A2(n223), .B1(ex_cp0_wdata[7]), 
        .B2(n283), .Z(n189) );
  AO22V4_8TH40 U80 ( .A1(mem_cp0_wdata[8]), .A2(n223), .B1(ex_cp0_wdata[8]), 
        .B2(n283), .Z(n190) );
  AO22V4_8TH40 U81 ( .A1(mem_cp0_wdata[9]), .A2(n223), .B1(ex_cp0_wdata[9]), 
        .B2(n283), .Z(n191) );
  AO22V4_8TH40 U82 ( .A1(mem_cp0_wdata[10]), .A2(n223), .B1(ex_cp0_wdata[10]), 
        .B2(n283), .Z(n192) );
  AO22V4_8TH40 U83 ( .A1(mem_cp0_wdata[11]), .A2(n223), .B1(ex_cp0_wdata[11]), 
        .B2(n283), .Z(n193) );
  AO22V4_8TH40 U84 ( .A1(mem_cp0_wdata[12]), .A2(n224), .B1(ex_cp0_wdata[12]), 
        .B2(n283), .Z(n194) );
  AO22V4_8TH40 U85 ( .A1(mem_cp0_wdata[13]), .A2(n224), .B1(ex_cp0_wdata[13]), 
        .B2(n283), .Z(n195) );
  AO22V4_8TH40 U86 ( .A1(mem_cp0_wdata[14]), .A2(n224), .B1(ex_cp0_wdata[14]), 
        .B2(n283), .Z(n196) );
  AO22V4_8TH40 U87 ( .A1(mem_cp0_wdata[15]), .A2(n224), .B1(ex_cp0_wdata[15]), 
        .B2(n283), .Z(n197) );
  AO22V4_8TH40 U88 ( .A1(mem_cp0_wdata[16]), .A2(n224), .B1(ex_cp0_wdata[16]), 
        .B2(n285), .Z(n198) );
  AO22V4_8TH40 U89 ( .A1(mem_cp0_wdata[17]), .A2(n224), .B1(ex_cp0_wdata[17]), 
        .B2(n288), .Z(n199) );
  AO22V4_8TH40 U90 ( .A1(mem_cp0_wdata[18]), .A2(n224), .B1(ex_cp0_wdata[18]), 
        .B2(n312), .Z(n200) );
  AO22V4_8TH40 U91 ( .A1(mem_cp0_wdata[19]), .A2(n224), .B1(ex_cp0_wdata[19]), 
        .B2(n247), .Z(n201) );
  AO22V4_8TH40 U92 ( .A1(mem_cp0_wdata[20]), .A2(n224), .B1(ex_cp0_wdata[20]), 
        .B2(n284), .Z(n202) );
  AO22V4_8TH40 U93 ( .A1(mem_cp0_wdata[21]), .A2(n224), .B1(ex_cp0_wdata[21]), 
        .B2(n290), .Z(n203) );
  AO22V4_8TH40 U94 ( .A1(mem_cp0_wdata[22]), .A2(n224), .B1(ex_cp0_wdata[22]), 
        .B2(n250), .Z(n204) );
  AO22V4_8TH40 U95 ( .A1(mem_cp0_wdata[23]), .A2(n224), .B1(ex_cp0_wdata[23]), 
        .B2(n286), .Z(n205) );
  AO22V4_8TH40 U96 ( .A1(mem_cp0_wdata[24]), .A2(n225), .B1(ex_cp0_wdata[24]), 
        .B2(n287), .Z(n206) );
  AO22V4_8TH40 U97 ( .A1(mem_cp0_wdata[25]), .A2(n225), .B1(ex_cp0_wdata[25]), 
        .B2(n289), .Z(n207) );
  AO22V4_8TH40 U98 ( .A1(mem_cp0_wdata[26]), .A2(n225), .B1(ex_cp0_wdata[26]), 
        .B2(n249), .Z(n208) );
  AO22V4_8TH40 U99 ( .A1(mem_cp0_wdata[27]), .A2(n225), .B1(ex_cp0_wdata[27]), 
        .B2(n284), .Z(n209) );
  AO22V4_8TH40 U100 ( .A1(mem_cp0_wdata[28]), .A2(n225), .B1(ex_cp0_wdata[28]), 
        .B2(n284), .Z(n210) );
  AO22V4_8TH40 U101 ( .A1(mem_cp0_wdata[29]), .A2(n225), .B1(ex_cp0_wdata[29]), 
        .B2(n284), .Z(n211) );
  AO22V4_8TH40 U102 ( .A1(mem_cp0_wdata[30]), .A2(n225), .B1(ex_cp0_wdata[30]), 
        .B2(n284), .Z(n212) );
  AO22V4_8TH40 U103 ( .A1(mem_cp0_wdata[31]), .A2(n225), .B1(ex_cp0_wdata[31]), 
        .B2(n284), .Z(n213) );
  AO22V4_8TH40 U104 ( .A1(mem_dmem_addr[31]), .A2(n235), .B1(ex_dmem_addr[31]), 
        .B2(n288), .Z(n69) );
  AO22V4_8TH40 U105 ( .A1(mem_dmem_addr[0]), .A2(n234), .B1(ex_dmem_addr[0]), 
        .B2(n287), .Z(n38) );
  AO22V4_8TH40 U106 ( .A1(mem_dmem_addr[1]), .A2(n234), .B1(ex_dmem_addr[1]), 
        .B2(n287), .Z(n39) );
  AO22V4_8TH40 U107 ( .A1(mem_dmem_addr[2]), .A2(n234), .B1(ex_dmem_addr[2]), 
        .B2(n287), .Z(n40) );
  AO22V4_8TH40 U108 ( .A1(mem_dmem_addr[3]), .A2(n234), .B1(ex_dmem_addr[3]), 
        .B2(n287), .Z(n41) );
  AO22V4_8TH40 U109 ( .A1(mem_dmem_addr[4]), .A2(n234), .B1(ex_dmem_addr[4]), 
        .B2(n287), .Z(n42) );
  AO22V4_8TH40 U110 ( .A1(mem_dmem_addr[5]), .A2(n234), .B1(ex_dmem_addr[5]), 
        .B2(n287), .Z(n43) );
  AO22V4_8TH40 U111 ( .A1(mem_dmem_addr[6]), .A2(n234), .B1(ex_dmem_addr[6]), 
        .B2(n287), .Z(n44) );
  AO22V4_8TH40 U112 ( .A1(mem_dmem_addr[7]), .A2(n234), .B1(ex_dmem_addr[7]), 
        .B2(n287), .Z(n45) );
  AO22V4_8TH40 U113 ( .A1(mem_dmem_addr[8]), .A2(n234), .B1(ex_dmem_addr[8]), 
        .B2(n283), .Z(n46) );
  AO22V4_8TH40 U114 ( .A1(mem_dmem_addr[9]), .A2(n234), .B1(ex_dmem_addr[9]), 
        .B2(n250), .Z(n47) );
  AO22V4_8TH40 U115 ( .A1(mem_dmem_addr[10]), .A2(n234), .B1(ex_dmem_addr[10]), 
        .B2(n285), .Z(n48) );
  AO22V4_8TH40 U116 ( .A1(mem_dmem_addr[11]), .A2(n219), .B1(ex_dmem_addr[11]), 
        .B2(n288), .Z(n49) );
  AO22V4_8TH40 U117 ( .A1(mem_dmem_addr[12]), .A2(n232), .B1(ex_dmem_addr[12]), 
        .B2(n312), .Z(n50) );
  AO22V4_8TH40 U118 ( .A1(mem_dmem_addr[13]), .A2(n220), .B1(ex_dmem_addr[13]), 
        .B2(n287), .Z(n51) );
  AO22V4_8TH40 U119 ( .A1(mem_dmem_addr[14]), .A2(n221), .B1(ex_dmem_addr[14]), 
        .B2(n248), .Z(n52) );
  AO22V4_8TH40 U120 ( .A1(mem_dmem_addr[15]), .A2(n224), .B1(ex_dmem_addr[15]), 
        .B2(n247), .Z(n53) );
  AO22V4_8TH40 U121 ( .A1(mem_dmem_addr[16]), .A2(n225), .B1(ex_dmem_addr[16]), 
        .B2(n284), .Z(n54) );
  AO22V4_8TH40 U122 ( .A1(mem_dmem_addr[17]), .A2(n236), .B1(ex_dmem_addr[17]), 
        .B2(n289), .Z(n55) );
  AO22V4_8TH40 U123 ( .A1(mem_dmem_addr[18]), .A2(n223), .B1(ex_dmem_addr[18]), 
        .B2(n290), .Z(n56) );
  AO22V4_8TH40 U124 ( .A1(mem_dmem_addr[19]), .A2(n3), .B1(ex_dmem_addr[19]), 
        .B2(n250), .Z(n57) );
  AO22V4_8TH40 U125 ( .A1(mem_dmem_addr[20]), .A2(n4), .B1(ex_dmem_addr[20]), 
        .B2(n285), .Z(n58) );
  AO22V4_8TH40 U126 ( .A1(mem_dmem_addr[21]), .A2(n235), .B1(ex_dmem_addr[21]), 
        .B2(n286), .Z(n59) );
  AO22V4_8TH40 U127 ( .A1(mem_dmem_addr[22]), .A2(n235), .B1(ex_dmem_addr[22]), 
        .B2(n288), .Z(n60) );
  AO22V4_8TH40 U128 ( .A1(mem_dmem_addr[23]), .A2(n235), .B1(ex_dmem_addr[23]), 
        .B2(n312), .Z(n61) );
  AO22V4_8TH40 U129 ( .A1(mem_dmem_addr[24]), .A2(n235), .B1(ex_dmem_addr[24]), 
        .B2(n287), .Z(n62) );
  AO22V4_8TH40 U130 ( .A1(mem_dmem_addr[25]), .A2(n235), .B1(ex_dmem_addr[25]), 
        .B2(n248), .Z(n63) );
  AO22V4_8TH40 U131 ( .A1(mem_dmem_addr[26]), .A2(n235), .B1(ex_dmem_addr[26]), 
        .B2(n247), .Z(n64) );
  AO22V4_8TH40 U132 ( .A1(mem_dmem_addr[27]), .A2(n235), .B1(ex_dmem_addr[27]), 
        .B2(n249), .Z(n65) );
  AO22V4_8TH40 U133 ( .A1(mem_dmem_addr[28]), .A2(n235), .B1(ex_dmem_addr[28]), 
        .B2(n284), .Z(n66) );
  AO22V4_8TH40 U134 ( .A1(mem_dmem_addr[29]), .A2(n235), .B1(ex_dmem_addr[29]), 
        .B2(n289), .Z(n67) );
  AO22V4_8TH40 U135 ( .A1(mem_dmem_addr[30]), .A2(n235), .B1(ex_dmem_addr[30]), 
        .B2(n288), .Z(n68) );
  AO22V4_8TH40 U136 ( .A1(mem_cp0_waddr[4]), .A2(n226), .B1(ex_cp0_waddr[4]), 
        .B2(n284), .Z(n218) );
  AO22V4_8TH40 U137 ( .A1(mem_cp0_waddr[3]), .A2(n225), .B1(ex_cp0_waddr[3]), 
        .B2(n284), .Z(n217) );
  AO22V4_8TH40 U138 ( .A1(mem_cp0_waddr[2]), .A2(n225), .B1(ex_cp0_waddr[2]), 
        .B2(n284), .Z(n216) );
  I2NOR3V2_8TH40 U139 ( .A1(flush_BAR), .A2(stall_ctrl[3]), .B(rst), .ZN(n313)
         );
  INV2_8TH40 U140 ( .I(n239), .ZN(n234) );
  INV2_8TH40 U141 ( .I(n238), .ZN(n235) );
  INV2_8TH40 U142 ( .I(n237), .ZN(n236) );
  INV2_8TH40 U143 ( .I(n246), .ZN(n2) );
  INV2_8TH40 U144 ( .I(n246), .ZN(n3) );
  INV2_8TH40 U145 ( .I(n245), .ZN(n4) );
  INV2_8TH40 U146 ( .I(n245), .ZN(n219) );
  INV2_8TH40 U147 ( .I(n244), .ZN(n220) );
  INV2_8TH40 U148 ( .I(n244), .ZN(n221) );
  INV2_8TH40 U149 ( .I(n243), .ZN(n222) );
  INV2_8TH40 U150 ( .I(n243), .ZN(n223) );
  INV2_8TH40 U151 ( .I(n242), .ZN(n224) );
  INV2_8TH40 U152 ( .I(n242), .ZN(n225) );
  INV2_8TH40 U153 ( .I(n241), .ZN(n226) );
  INV2_8TH40 U154 ( .I(n240), .ZN(n232) );
  INV2_8TH40 U155 ( .I(n240), .ZN(n233) );
  CLKBUFV2_8TH40 U156 ( .I(n1), .Z(n239) );
  CLKBUFV2_8TH40 U157 ( .I(n242), .Z(n238) );
  CLKBUFV2_8TH40 U158 ( .I(n241), .Z(n237) );
  CLKBUFV2_8TH40 U159 ( .I(n240), .Z(n242) );
  CLKBUFV2_8TH40 U160 ( .I(n243), .Z(n241) );
  CLKBUFV2_8TH40 U161 ( .I(n244), .Z(n240) );
  CLKBUFV2_8TH40 U162 ( .I(n245), .Z(n246) );
  CLKBUFV2_8TH40 U163 ( .I(n239), .Z(n245) );
  CLKBUFV2_8TH40 U164 ( .I(n1), .Z(n244) );
  CLKBUFV2_8TH40 U165 ( .I(n1), .Z(n243) );
  INV2_8TH40 U166 ( .I(n293), .ZN(n287) );
  INV2_8TH40 U167 ( .I(n292), .ZN(n288) );
  INV2_8TH40 U168 ( .I(n300), .ZN(n248) );
  INV2_8TH40 U169 ( .I(n299), .ZN(n249) );
  INV2_8TH40 U170 ( .I(n298), .ZN(n250) );
  INV2_8TH40 U171 ( .I(n297), .ZN(n283) );
  INV2_8TH40 U172 ( .I(n296), .ZN(n284) );
  INV2_8TH40 U173 ( .I(n295), .ZN(n285) );
  INV2_8TH40 U174 ( .I(n294), .ZN(n286) );
  CLKBUFV2_8TH40 U175 ( .I(n306), .Z(n293) );
  CLKBUFV2_8TH40 U176 ( .I(n306), .Z(n292) );
  CLKBUFV2_8TH40 U177 ( .I(n302), .Z(n300) );
  CLKBUFV2_8TH40 U178 ( .I(n303), .Z(n299) );
  CLKBUFV2_8TH40 U179 ( .I(n303), .Z(n298) );
  CLKBUFV2_8TH40 U180 ( .I(n304), .Z(n297) );
  CLKBUFV2_8TH40 U181 ( .I(n304), .Z(n296) );
  CLKBUFV2_8TH40 U182 ( .I(n305), .Z(n295) );
  CLKBUFV2_8TH40 U183 ( .I(n305), .Z(n294) );
  INV2_8TH40 U184 ( .I(n291), .ZN(n289) );
  INV2_8TH40 U185 ( .I(n291), .ZN(n290) );
  INV2_8TH40 U186 ( .I(n301), .ZN(n247) );
  CLKBUFV2_8TH40 U187 ( .I(n302), .Z(n301) );
  BUFV4_8TH40 U188 ( .I(n307), .Z(n291) );
  CLKBUFV2_8TH40 U189 ( .I(n308), .Z(n307) );
  CLKBUFV2_8TH40 U190 ( .I(n308), .Z(n306) );
  CLKBUFV2_8TH40 U191 ( .I(n310), .Z(n302) );
  CLKBUFV2_8TH40 U192 ( .I(n310), .Z(n303) );
  CLKBUFV2_8TH40 U193 ( .I(n309), .Z(n304) );
  CLKBUFV2_8TH40 U194 ( .I(n309), .Z(n305) );
  CLKBUFV2_8TH40 U195 ( .I(n311), .Z(n308) );
  CLKBUFV2_8TH40 U196 ( .I(n311), .Z(n310) );
  CLKBUFV2_8TH40 U197 ( .I(n311), .Z(n309) );
  INV2_8TH40 U198 ( .I(n312), .ZN(n311) );
  AO22V0_8TH40 U199 ( .A1(mem_ls_data_tmp[3]), .A2(n236), .B1(
        ex_ls_data_tmp[3]), .B2(n290), .Z(n9) );
  AO22V0_8TH40 U200 ( .A1(mem_ls_data_tmp[2]), .A2(n233), .B1(
        ex_ls_data_tmp[2]), .B2(n289), .Z(n8) );
  AO22V0_8TH40 U201 ( .A1(mem_inst_type[7]), .A2(n235), .B1(ex_inst_type[7]), 
        .B2(n288), .Z(n77) );
  AO22V0_8TH40 U202 ( .A1(mem_inst_type[6]), .A2(n226), .B1(ex_inst_type[6]), 
        .B2(n288), .Z(n76) );
  AO22V0_8TH40 U203 ( .A1(mem_inst_type[5]), .A2(n222), .B1(ex_inst_type[5]), 
        .B2(n288), .Z(n75) );
  AO22V0_8TH40 U204 ( .A1(mem_inst_type[4]), .A2(n233), .B1(ex_inst_type[4]), 
        .B2(n288), .Z(n74) );
  AO22V0_8TH40 U205 ( .A1(mem_inst_type[3]), .A2(n2), .B1(ex_inst_type[3]), 
        .B2(n288), .Z(n73) );
  AO22V0_8TH40 U206 ( .A1(mem_inst_type[2]), .A2(n234), .B1(ex_inst_type[2]), 
        .B2(n288), .Z(n72) );
  AO22V0_8TH40 U207 ( .A1(mem_inst_type[1]), .A2(n235), .B1(ex_inst_type[1]), 
        .B2(n288), .Z(n71) );
  AO22V0_8TH40 U208 ( .A1(mem_inst_type[0]), .A2(n235), .B1(ex_inst_type[0]), 
        .B2(n288), .Z(n70) );
  AO22V0_8TH40 U209 ( .A1(mem_ls_data_tmp[1]), .A2(n235), .B1(
        ex_ls_data_tmp[1]), .B2(n288), .Z(n7) );
  AO22V0_8TH40 U210 ( .A1(mem_ls_data_tmp[0]), .A2(n226), .B1(
        ex_ls_data_tmp[0]), .B2(n285), .Z(n6) );
  AO22V0_8TH40 U211 ( .A1(mem_cp0_we), .A2(n233), .B1(ex_cp0_we), .B2(n249), 
        .Z(n5) );
  AO22V0_8TH40 U212 ( .A1(mem_ls_data_tmp[31]), .A2(n234), .B1(
        ex_ls_data_tmp[31]), .B2(n287), .Z(n37) );
  AO22V0_8TH40 U213 ( .A1(mem_ls_data_tmp[30]), .A2(n234), .B1(
        ex_ls_data_tmp[30]), .B2(n287), .Z(n36) );
  AO22V0_8TH40 U214 ( .A1(mem_ls_data_tmp[29]), .A2(n233), .B1(
        ex_ls_data_tmp[29]), .B2(n287), .Z(n35) );
  AO22V0_8TH40 U215 ( .A1(mem_ls_data_tmp[28]), .A2(n233), .B1(
        ex_ls_data_tmp[28]), .B2(n287), .Z(n34) );
  AO22V0_8TH40 U216 ( .A1(mem_ls_data_tmp[27]), .A2(n233), .B1(
        ex_ls_data_tmp[27]), .B2(n286), .Z(n33) );
  AO22V0_8TH40 U217 ( .A1(mem_ls_data_tmp[26]), .A2(n233), .B1(
        ex_ls_data_tmp[26]), .B2(n286), .Z(n32) );
  AO22V0_8TH40 U218 ( .A1(mem_ls_data_tmp[25]), .A2(n233), .B1(
        ex_ls_data_tmp[25]), .B2(n286), .Z(n31) );
  AO22V0_8TH40 U219 ( .A1(mem_ls_data_tmp[24]), .A2(n233), .B1(
        ex_ls_data_tmp[24]), .B2(n286), .Z(n30) );
  AO22V0_8TH40 U220 ( .A1(mem_ls_data_tmp[23]), .A2(n233), .B1(
        ex_ls_data_tmp[23]), .B2(n286), .Z(n29) );
  AO22V0_8TH40 U221 ( .A1(mem_cur_inst_addr[31]), .A2(n233), .B1(
        ex_cur_inst_addr[31]), .B2(n286), .Z(n282) );
  AO22V0_8TH40 U222 ( .A1(mem_cur_inst_addr[30]), .A2(n233), .B1(
        ex_cur_inst_addr[30]), .B2(n286), .Z(n281) );
  AO22V0_8TH40 U223 ( .A1(mem_cur_inst_addr[29]), .A2(n233), .B1(
        ex_cur_inst_addr[29]), .B2(n286), .Z(n280) );
  AO22V0_8TH40 U224 ( .A1(mem_ls_data_tmp[22]), .A2(n233), .B1(
        ex_ls_data_tmp[22]), .B2(n286), .Z(n28) );
  AO22V0_8TH40 U225 ( .A1(mem_cur_inst_addr[28]), .A2(n233), .B1(
        ex_cur_inst_addr[28]), .B2(n286), .Z(n279) );
  AO22V0_8TH40 U226 ( .A1(mem_cur_inst_addr[27]), .A2(n233), .B1(
        ex_cur_inst_addr[27]), .B2(n286), .Z(n278) );
  AO22V0_8TH40 U227 ( .A1(mem_cur_inst_addr[26]), .A2(n232), .B1(
        ex_cur_inst_addr[26]), .B2(n286), .Z(n277) );
  AO22V0_8TH40 U228 ( .A1(mem_cur_inst_addr[25]), .A2(n232), .B1(
        ex_cur_inst_addr[25]), .B2(n247), .Z(n276) );
  AO22V0_8TH40 U229 ( .A1(mem_cur_inst_addr[24]), .A2(n232), .B1(
        ex_cur_inst_addr[24]), .B2(n284), .Z(n275) );
  AO22V0_8TH40 U230 ( .A1(mem_cur_inst_addr[23]), .A2(n232), .B1(
        ex_cur_inst_addr[23]), .B2(n290), .Z(n274) );
  AO22V0_8TH40 U231 ( .A1(mem_cur_inst_addr[22]), .A2(n232), .B1(
        ex_cur_inst_addr[22]), .B2(n287), .Z(n273) );
  AO22V0_8TH40 U232 ( .A1(mem_cur_inst_addr[21]), .A2(n232), .B1(
        ex_cur_inst_addr[21]), .B2(n289), .Z(n272) );
  AO22V0_8TH40 U233 ( .A1(mem_cur_inst_addr[20]), .A2(n232), .B1(
        ex_cur_inst_addr[20]), .B2(n286), .Z(n271) );
  AO22V0_8TH40 U234 ( .A1(mem_cur_inst_addr[19]), .A2(n232), .B1(
        ex_cur_inst_addr[19]), .B2(n250), .Z(n270) );
  AO22V0_8TH40 U235 ( .A1(mem_ls_data_tmp[21]), .A2(n232), .B1(
        ex_ls_data_tmp[21]), .B2(n248), .Z(n27) );
  AO22V0_8TH40 U236 ( .A1(mem_cur_inst_addr[18]), .A2(n232), .B1(
        ex_cur_inst_addr[18]), .B2(n287), .Z(n269) );
  AO22V0_8TH40 U237 ( .A1(mem_cur_inst_addr[17]), .A2(n232), .B1(
        ex_cur_inst_addr[17]), .B2(n249), .Z(n268) );
  AO22V0_8TH40 U238 ( .A1(mem_cur_inst_addr[16]), .A2(n232), .B1(
        ex_cur_inst_addr[16]), .B2(n283), .Z(n267) );
  AO22V0_8TH40 U239 ( .A1(mem_cur_inst_addr[15]), .A2(n232), .B1(
        ex_cur_inst_addr[15]), .B2(n283), .Z(n266) );
  AO22V0_8TH40 U240 ( .A1(mem_cur_inst_addr[14]), .A2(n222), .B1(
        ex_cur_inst_addr[14]), .B2(n285), .Z(n265) );
  AO22V0_8TH40 U241 ( .A1(mem_cur_inst_addr[13]), .A2(n226), .B1(
        ex_cur_inst_addr[13]), .B2(n285), .Z(n264) );
  AO22V0_8TH40 U242 ( .A1(mem_cur_inst_addr[12]), .A2(n222), .B1(
        ex_cur_inst_addr[12]), .B2(n285), .Z(n263) );
  AO22V0_8TH40 U243 ( .A1(mem_cur_inst_addr[11]), .A2(n232), .B1(
        ex_cur_inst_addr[11]), .B2(n285), .Z(n262) );
  AO22V0_8TH40 U244 ( .A1(mem_cur_inst_addr[10]), .A2(n233), .B1(
        ex_cur_inst_addr[10]), .B2(n285), .Z(n261) );
  AO22V0_8TH40 U245 ( .A1(mem_cur_inst_addr[9]), .A2(n220), .B1(
        ex_cur_inst_addr[9]), .B2(n285), .Z(n260) );
  AO22V0_8TH40 U246 ( .A1(mem_ls_data_tmp[20]), .A2(n221), .B1(
        ex_ls_data_tmp[20]), .B2(n285), .Z(n26) );
  AO22V0_8TH40 U247 ( .A1(mem_cur_inst_addr[8]), .A2(n226), .B1(
        ex_cur_inst_addr[8]), .B2(n285), .Z(n259) );
  AO22V0_8TH40 U248 ( .A1(mem_cur_inst_addr[7]), .A2(n222), .B1(
        ex_cur_inst_addr[7]), .B2(n285), .Z(n258) );
  AO22V0_8TH40 U249 ( .A1(mem_cur_inst_addr[6]), .A2(n232), .B1(
        ex_cur_inst_addr[6]), .B2(n285), .Z(n257) );
  AO22V0_8TH40 U250 ( .A1(mem_cur_inst_addr[5]), .A2(n233), .B1(
        ex_cur_inst_addr[5]), .B2(n285), .Z(n256) );
  AO22V0_8TH40 U251 ( .A1(mem_cur_inst_addr[4]), .A2(n220), .B1(
        ex_cur_inst_addr[4]), .B2(n285), .Z(n255) );
  AO22V0_8TH40 U252 ( .A1(mem_cur_inst_addr[3]), .A2(n221), .B1(
        ex_cur_inst_addr[3]), .B2(n284), .Z(n254) );
  AO22V0_8TH40 U253 ( .A1(mem_cur_inst_addr[2]), .A2(n226), .B1(
        ex_cur_inst_addr[2]), .B2(n290), .Z(n253) );
  AO22V0_8TH40 U254 ( .A1(mem_cur_inst_addr[1]), .A2(n226), .B1(
        ex_cur_inst_addr[1]), .B2(n286), .Z(n252) );
  AO22V0_8TH40 U255 ( .A1(mem_cur_inst_addr[0]), .A2(n226), .B1(
        ex_cur_inst_addr[0]), .B2(n287), .Z(n251) );
  AO22V0_8TH40 U256 ( .A1(mem_ls_data_tmp[19]), .A2(n226), .B1(
        ex_ls_data_tmp[19]), .B2(n289), .Z(n25) );
  AO22V0_8TH40 U257 ( .A1(mem_ls_data_tmp[18]), .A2(n226), .B1(
        ex_ls_data_tmp[18]), .B2(n290), .Z(n24) );
  AO22V0_8TH40 U258 ( .A1(mem_except_type[12]), .A2(n226), .B1(
        ex_except_type[12]), .B2(n290), .Z(n231) );
  AO22V0_8TH40 U259 ( .A1(mem_except_type[11]), .A2(n226), .B1(
        ex_except_type[11]), .B2(n248), .Z(n230) );
  AO22V0_8TH40 U260 ( .A1(mem_ls_data_tmp[17]), .A2(n226), .B1(
        ex_ls_data_tmp[17]), .B2(n250), .Z(n23) );
  AO22V0_8TH40 U261 ( .A1(mem_except_type[9]), .A2(n226), .B1(
        ex_except_type[9]), .B2(n249), .Z(n228) );
  AO22V0_8TH40 U262 ( .A1(mem_except_type[8]), .A2(n226), .B1(
        ex_except_type[8]), .B2(n283), .Z(n227) );
  AO22V0_8TH40 U263 ( .A1(mem_ls_data_tmp[16]), .A2(n226), .B1(
        ex_ls_data_tmp[16]), .B2(n284), .Z(n22) );
  AO22V0_8TH40 U264 ( .A1(mem_ls_data_tmp[15]), .A2(n225), .B1(
        ex_ls_data_tmp[15]), .B2(n284), .Z(n21) );
  AO22V0_8TH40 U265 ( .A1(mem_ls_data_tmp[14]), .A2(n224), .B1(
        ex_ls_data_tmp[14]), .B2(n248), .Z(n20) );
  AO22V0_8TH40 U266 ( .A1(mem_ls_data_tmp[13]), .A2(n223), .B1(
        ex_ls_data_tmp[13]), .B2(n283), .Z(n19) );
  AO22V0_8TH40 U267 ( .A1(mem_inst_delayslot), .A2(n222), .B1(
        ex_inst_delayslot), .B2(n285), .Z(n181) );
  AO22V0_8TH40 U268 ( .A1(mem_gpr_we), .A2(n222), .B1(ex_gpr_we), .B2(n312), 
        .Z(n180) );
  AO22V0_8TH40 U269 ( .A1(mem_ls_data_tmp[12]), .A2(n222), .B1(
        ex_ls_data_tmp[12]), .B2(n290), .Z(n18) );
  AO22V0_8TH40 U270 ( .A1(mem_target_gpr[4]), .A2(n222), .B1(ex_target_gpr[4]), 
        .B2(n287), .Z(n179) );
  AO22V0_8TH40 U271 ( .A1(mem_target_gpr[3]), .A2(n222), .B1(ex_target_gpr[3]), 
        .B2(n250), .Z(n178) );
  AO22V0_8TH40 U272 ( .A1(mem_target_gpr[2]), .A2(n222), .B1(ex_target_gpr[2]), 
        .B2(n288), .Z(n177) );
  AO22V0_8TH40 U273 ( .A1(mem_target_gpr[1]), .A2(n222), .B1(ex_target_gpr[1]), 
        .B2(n285), .Z(n176) );
  AO22V0_8TH40 U274 ( .A1(mem_target_gpr[0]), .A2(n222), .B1(ex_target_gpr[0]), 
        .B2(n250), .Z(n175) );
  AO22V0_8TH40 U275 ( .A1(mem_exe_result[31]), .A2(n222), .B1(
        ex_exe_result[31]), .B2(n250), .Z(n174) );
  AO22V0_8TH40 U276 ( .A1(mem_exe_result[30]), .A2(n222), .B1(
        ex_exe_result[30]), .B2(n250), .Z(n173) );
  AO22V0_8TH40 U277 ( .A1(mem_exe_result[29]), .A2(n222), .B1(
        ex_exe_result[29]), .B2(n250), .Z(n172) );
  AO22V0_8TH40 U278 ( .A1(mem_exe_result[28]), .A2(n222), .B1(
        ex_exe_result[28]), .B2(n250), .Z(n171) );
  AO22V0_8TH40 U279 ( .A1(mem_exe_result[27]), .A2(n222), .B1(
        ex_exe_result[27]), .B2(n250), .Z(n170) );
  AO22V0_8TH40 U280 ( .A1(mem_ls_data_tmp[11]), .A2(n221), .B1(
        ex_ls_data_tmp[11]), .B2(n250), .Z(n17) );
  AO22V0_8TH40 U281 ( .A1(mem_exe_result[26]), .A2(n221), .B1(
        ex_exe_result[26]), .B2(n250), .Z(n169) );
  AO22V0_8TH40 U282 ( .A1(mem_exe_result[25]), .A2(n221), .B1(
        ex_exe_result[25]), .B2(n250), .Z(n168) );
  AO22V0_8TH40 U283 ( .A1(mem_exe_result[24]), .A2(n221), .B1(
        ex_exe_result[24]), .B2(n250), .Z(n167) );
  AO22V0_8TH40 U284 ( .A1(mem_exe_result[23]), .A2(n221), .B1(
        ex_exe_result[23]), .B2(n250), .Z(n166) );
  AO22V0_8TH40 U285 ( .A1(mem_exe_result[22]), .A2(n221), .B1(
        ex_exe_result[22]), .B2(n250), .Z(n165) );
  AO22V0_8TH40 U286 ( .A1(mem_exe_result[21]), .A2(n221), .B1(
        ex_exe_result[21]), .B2(n288), .Z(n164) );
  AO22V0_8TH40 U287 ( .A1(mem_exe_result[20]), .A2(n221), .B1(
        ex_exe_result[20]), .B2(n286), .Z(n163) );
  AO22V0_8TH40 U288 ( .A1(mem_exe_result[19]), .A2(n221), .B1(
        ex_exe_result[19]), .B2(n250), .Z(n162) );
  AO22V0_8TH40 U289 ( .A1(mem_exe_result[18]), .A2(n221), .B1(
        ex_exe_result[18]), .B2(n312), .Z(n161) );
  AO22V0_8TH40 U290 ( .A1(mem_exe_result[17]), .A2(n221), .B1(
        ex_exe_result[17]), .B2(n312), .Z(n160) );
  AO22V0_8TH40 U291 ( .A1(mem_ls_data_tmp[10]), .A2(n221), .B1(
        ex_ls_data_tmp[10]), .B2(n285), .Z(n16) );
  AO22V0_8TH40 U292 ( .A1(mem_exe_result[16]), .A2(n221), .B1(
        ex_exe_result[16]), .B2(n312), .Z(n159) );
  AO22V0_8TH40 U293 ( .A1(mem_exe_result[15]), .A2(n220), .B1(
        ex_exe_result[15]), .B2(n286), .Z(n158) );
  AO22V0_8TH40 U294 ( .A1(mem_exe_result[14]), .A2(n220), .B1(
        ex_exe_result[14]), .B2(n250), .Z(n157) );
  AO22V0_8TH40 U295 ( .A1(mem_exe_result[13]), .A2(n220), .B1(
        ex_exe_result[13]), .B2(n288), .Z(n156) );
  AO22V0_8TH40 U296 ( .A1(mem_exe_result[12]), .A2(n220), .B1(
        ex_exe_result[12]), .B2(n247), .Z(n155) );
  AO22V0_8TH40 U297 ( .A1(mem_exe_result[11]), .A2(n220), .B1(
        ex_exe_result[11]), .B2(n312), .Z(n154) );
  AO22V0_8TH40 U298 ( .A1(mem_exe_result[10]), .A2(n220), .B1(
        ex_exe_result[10]), .B2(n312), .Z(n153) );
  AO22V0_8TH40 U299 ( .A1(mem_exe_result[9]), .A2(n220), .B1(ex_exe_result[9]), 
        .B2(n312), .Z(n152) );
  AO22V0_8TH40 U300 ( .A1(mem_exe_result[8]), .A2(n220), .B1(ex_exe_result[8]), 
        .B2(n312), .Z(n151) );
  AO22V0_8TH40 U301 ( .A1(mem_exe_result[7]), .A2(n220), .B1(ex_exe_result[7]), 
        .B2(n312), .Z(n150) );
  AO22V0_8TH40 U302 ( .A1(mem_ls_data_tmp[9]), .A2(n220), .B1(
        ex_ls_data_tmp[9]), .B2(n312), .Z(n15) );
  AO22V0_8TH40 U303 ( .A1(mem_exe_result[6]), .A2(n220), .B1(ex_exe_result[6]), 
        .B2(n312), .Z(n149) );
  AO22V0_8TH40 U304 ( .A1(mem_exe_result[5]), .A2(n220), .B1(ex_exe_result[5]), 
        .B2(n312), .Z(n148) );
  AO22V0_8TH40 U305 ( .A1(mem_exe_result[4]), .A2(n220), .B1(ex_exe_result[4]), 
        .B2(n312), .Z(n147) );
  AO22V0_8TH40 U306 ( .A1(mem_exe_result[3]), .A2(n219), .B1(ex_exe_result[3]), 
        .B2(n312), .Z(n146) );
  AO22V0_8TH40 U307 ( .A1(mem_exe_result[2]), .A2(n219), .B1(ex_exe_result[2]), 
        .B2(n312), .Z(n145) );
  AO22V0_8TH40 U308 ( .A1(mem_exe_result[1]), .A2(n219), .B1(ex_exe_result[1]), 
        .B2(n312), .Z(n144) );
  AO22V0_8TH40 U309 ( .A1(mem_exe_result[0]), .A2(n219), .B1(ex_exe_result[0]), 
        .B2(n285), .Z(n143) );
  AO22V0_8TH40 U310 ( .A1(mem_ls_data_tmp[8]), .A2(n219), .B1(
        ex_ls_data_tmp[8]), .B2(n249), .Z(n14) );
  AO22V0_8TH40 U311 ( .A1(mem_ls_data_tmp[7]), .A2(n4), .B1(ex_ls_data_tmp[7]), 
        .B2(n289), .Z(n13) );
  AO22V0_8TH40 U312 ( .A1(mem_ls_data_tmp[6]), .A2(n3), .B1(ex_ls_data_tmp[6]), 
        .B2(n248), .Z(n12) );
  AO22V0_8TH40 U313 ( .A1(mem_ls_data_tmp[5]), .A2(n2), .B1(ex_ls_data_tmp[5]), 
        .B2(n247), .Z(n11) );
  AO22V0_8TH40 U314 ( .A1(mem_ls_data_tmp[4]), .A2(n2), .B1(ex_ls_data_tmp[4]), 
        .B2(n247), .Z(n10) );
  INOR3V0_8TH40 U315 ( .A1(flush_BAR), .B1(rst), .B2(stall_ctrl[3]), .ZN(n312)
         );
endmodule


module mem_access ( rst, gpr_we, target_gpr, exe_result, hi, lo, hilo_we, 
        inst_type, ls_data_tmp, dmem_addr_i, dmem_data_i, llbit_i, wb_llbit_we, 
        wb_llbit_value, cp0_we_i, cp0_waddr_i, cp0_wdata_i, except_type_i, 
        in_delayslot_i, cur_inst_addr_i, cp0_status_i, cp0_cause_i, cp0_epc_i, 
        wb_cp0_we, wb_cp0_waddr, wb_cp0_wdata, dmem_addr_o, dmem_data_o, 
        dmem_byte_sel, dmem_ce, dmem_we, gpr_we_o, target_gpr_o, exe_result_o, 
        hi_o, lo_o, hilo_we_o, mem_llbit_we, mem_llbit_value, cp0_we_o, 
        cp0_waddr_o, cp0_wdata_o, except_type_o, cp0_epc_o, cur_inst_addr_o, 
        in_delayslot_o );
  input [4:0] target_gpr;
  input [31:0] exe_result;
  input [31:0] hi;
  input [31:0] lo;
  input [7:0] inst_type;
  input [31:0] ls_data_tmp;
  input [31:0] dmem_addr_i;
  input [31:0] dmem_data_i;
  input [4:0] cp0_waddr_i;
  input [31:0] cp0_wdata_i;
  input [31:0] except_type_i;
  input [31:0] cur_inst_addr_i;
  input [31:0] cp0_status_i;
  input [31:0] cp0_cause_i;
  input [31:0] cp0_epc_i;
  input [4:0] wb_cp0_waddr;
  input [31:0] wb_cp0_wdata;
  output [31:0] dmem_addr_o;
  output [31:0] dmem_data_o;
  output [3:0] dmem_byte_sel;
  output [4:0] target_gpr_o;
  output [31:0] exe_result_o;
  output [31:0] hi_o;
  output [31:0] lo_o;
  output [4:0] cp0_waddr_o;
  output [31:0] cp0_wdata_o;
  output [31:0] except_type_o;
  output [31:0] cp0_epc_o;
  output [31:0] cur_inst_addr_o;
  input rst, gpr_we, hilo_we, llbit_i, wb_llbit_we, wb_llbit_value, cp0_we_i,
         in_delayslot_i, wb_cp0_we;
  output dmem_ce, dmem_we, gpr_we_o, hilo_we_o, mem_llbit_we, mem_llbit_value,
         cp0_we_o, in_delayslot_o;
  wire   in_delayslot_i, N569, N570, N571, N572, N573, N574, N575, N576, N577,
         N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588,
         N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599,
         N600, N601, n333, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352;
  wire   [15:10] cp0_cause;
  assign cur_inst_addr_o[31] = cur_inst_addr_i[31];
  assign cur_inst_addr_o[30] = cur_inst_addr_i[30];
  assign cur_inst_addr_o[29] = cur_inst_addr_i[29];
  assign cur_inst_addr_o[28] = cur_inst_addr_i[28];
  assign cur_inst_addr_o[27] = cur_inst_addr_i[27];
  assign cur_inst_addr_o[26] = cur_inst_addr_i[26];
  assign cur_inst_addr_o[25] = cur_inst_addr_i[25];
  assign cur_inst_addr_o[24] = cur_inst_addr_i[24];
  assign cur_inst_addr_o[23] = cur_inst_addr_i[23];
  assign cur_inst_addr_o[22] = cur_inst_addr_i[22];
  assign cur_inst_addr_o[21] = cur_inst_addr_i[21];
  assign cur_inst_addr_o[20] = cur_inst_addr_i[20];
  assign cur_inst_addr_o[19] = cur_inst_addr_i[19];
  assign cur_inst_addr_o[18] = cur_inst_addr_i[18];
  assign cur_inst_addr_o[17] = cur_inst_addr_i[17];
  assign cur_inst_addr_o[16] = cur_inst_addr_i[16];
  assign cur_inst_addr_o[15] = cur_inst_addr_i[15];
  assign cur_inst_addr_o[14] = cur_inst_addr_i[14];
  assign cur_inst_addr_o[13] = cur_inst_addr_i[13];
  assign cur_inst_addr_o[12] = cur_inst_addr_i[12];
  assign cur_inst_addr_o[11] = cur_inst_addr_i[11];
  assign cur_inst_addr_o[10] = cur_inst_addr_i[10];
  assign cur_inst_addr_o[9] = cur_inst_addr_i[9];
  assign cur_inst_addr_o[8] = cur_inst_addr_i[8];
  assign cur_inst_addr_o[7] = cur_inst_addr_i[7];
  assign cur_inst_addr_o[6] = cur_inst_addr_i[6];
  assign cur_inst_addr_o[5] = cur_inst_addr_i[5];
  assign cur_inst_addr_o[4] = cur_inst_addr_i[4];
  assign cur_inst_addr_o[3] = cur_inst_addr_i[3];
  assign cur_inst_addr_o[2] = cur_inst_addr_i[2];
  assign cur_inst_addr_o[1] = cur_inst_addr_i[1];
  assign cur_inst_addr_o[0] = cur_inst_addr_i[0];
  assign in_delayslot_o = in_delayslot_i;

  LAHRNQV1_8TH40 cp0_cause_reg_15_ ( .E(n333), .D(cp0_cause_i[15]), .RDN(n352), 
        .Q(cp0_cause[15]) );
  LAHRNQV1_8TH40 cp0_cause_reg_14_ ( .E(n333), .D(cp0_cause_i[14]), .RDN(n352), 
        .Q(cp0_cause[14]) );
  LAHRNQV1_8TH40 cp0_cause_reg_13_ ( .E(n333), .D(cp0_cause_i[13]), .RDN(n352), 
        .Q(cp0_cause[13]) );
  LAHRNQV1_8TH40 cp0_cause_reg_12_ ( .E(n333), .D(cp0_cause_i[12]), .RDN(n352), 
        .Q(cp0_cause[12]) );
  LAHRNQV1_8TH40 cp0_cause_reg_11_ ( .E(n333), .D(cp0_cause_i[11]), .RDN(n352), 
        .Q(cp0_cause[11]) );
  LAHRNQV1_8TH40 cp0_cause_reg_10_ ( .E(n333), .D(cp0_cause_i[10]), .RDN(n352), 
        .Q(cp0_cause[10]) );
  LAHQV4_8TH40 dmem_data_o_reg_31_ ( .E(N569), .D(N601), .Q(dmem_data_o[31])
         );
  LAHQV4_8TH40 dmem_data_o_reg_30_ ( .E(N569), .D(N600), .Q(dmem_data_o[30])
         );
  LAHQV4_8TH40 dmem_data_o_reg_29_ ( .E(N569), .D(N599), .Q(dmem_data_o[29])
         );
  LAHQV4_8TH40 dmem_data_o_reg_28_ ( .E(N569), .D(N598), .Q(dmem_data_o[28])
         );
  LAHQV4_8TH40 dmem_data_o_reg_27_ ( .E(N569), .D(N597), .Q(dmem_data_o[27])
         );
  LAHQV4_8TH40 dmem_data_o_reg_26_ ( .E(N569), .D(N596), .Q(dmem_data_o[26])
         );
  LAHQV4_8TH40 dmem_data_o_reg_25_ ( .E(N569), .D(N595), .Q(dmem_data_o[25])
         );
  LAHQV4_8TH40 dmem_data_o_reg_24_ ( .E(N569), .D(N594), .Q(dmem_data_o[24])
         );
  LAHQV4_8TH40 dmem_data_o_reg_23_ ( .E(N569), .D(N593), .Q(dmem_data_o[23])
         );
  LAHQV4_8TH40 dmem_data_o_reg_22_ ( .E(N569), .D(N592), .Q(dmem_data_o[22])
         );
  LAHQV4_8TH40 dmem_data_o_reg_21_ ( .E(N569), .D(N591), .Q(dmem_data_o[21])
         );
  LAHQV4_8TH40 dmem_data_o_reg_20_ ( .E(N569), .D(N590), .Q(dmem_data_o[20])
         );
  LAHQV4_8TH40 dmem_data_o_reg_19_ ( .E(N569), .D(N589), .Q(dmem_data_o[19])
         );
  LAHQV4_8TH40 dmem_data_o_reg_18_ ( .E(N569), .D(N588), .Q(dmem_data_o[18])
         );
  LAHQV4_8TH40 dmem_data_o_reg_17_ ( .E(N569), .D(N587), .Q(dmem_data_o[17])
         );
  LAHQV4_8TH40 dmem_data_o_reg_16_ ( .E(N569), .D(N586), .Q(dmem_data_o[16])
         );
  LAHQV4_8TH40 dmem_data_o_reg_15_ ( .E(N569), .D(N585), .Q(dmem_data_o[15])
         );
  LAHQV4_8TH40 dmem_data_o_reg_14_ ( .E(N569), .D(N584), .Q(dmem_data_o[14])
         );
  LAHQV4_8TH40 dmem_data_o_reg_13_ ( .E(N569), .D(N583), .Q(dmem_data_o[13])
         );
  LAHQV4_8TH40 dmem_data_o_reg_12_ ( .E(N569), .D(N582), .Q(dmem_data_o[12])
         );
  LAHQV4_8TH40 dmem_data_o_reg_11_ ( .E(N569), .D(N581), .Q(dmem_data_o[11])
         );
  LAHQV4_8TH40 dmem_data_o_reg_10_ ( .E(N569), .D(N580), .Q(dmem_data_o[10])
         );
  LAHQV4_8TH40 dmem_data_o_reg_9_ ( .E(N569), .D(N579), .Q(dmem_data_o[9]) );
  LAHQV4_8TH40 dmem_data_o_reg_8_ ( .E(N569), .D(N578), .Q(dmem_data_o[8]) );
  LAHQV4_8TH40 dmem_data_o_reg_7_ ( .E(N569), .D(N577), .Q(dmem_data_o[7]) );
  LAHQV4_8TH40 dmem_data_o_reg_6_ ( .E(N569), .D(N576), .Q(dmem_data_o[6]) );
  LAHQV4_8TH40 dmem_data_o_reg_5_ ( .E(N569), .D(N575), .Q(dmem_data_o[5]) );
  LAHQV4_8TH40 dmem_data_o_reg_4_ ( .E(N569), .D(N574), .Q(dmem_data_o[4]) );
  LAHQV4_8TH40 dmem_data_o_reg_3_ ( .E(N569), .D(N573), .Q(dmem_data_o[3]) );
  LAHQV4_8TH40 dmem_data_o_reg_2_ ( .E(N569), .D(N572), .Q(dmem_data_o[2]) );
  LAHQV4_8TH40 dmem_data_o_reg_1_ ( .E(N569), .D(N571), .Q(dmem_data_o[1]) );
  LAHQV4_8TH40 dmem_data_o_reg_0_ ( .E(N569), .D(N570), .Q(dmem_data_o[0]) );
  AO221V4_8TH40 U3 ( .A1(n252), .A2(n256), .B1(n352), .B2(n259), .C(n260), .Z(
        dmem_byte_sel[0]) );
  AND2V4_8TH40 U4 ( .A1(n229), .A2(n230), .Z(n225) );
  NAND3V2_8TH40 U5 ( .A1(n271), .A2(n65), .A3(n272), .ZN(dmem_ce) );
  OAI21V2_8TH40 U6 ( .A1(n201), .A2(n4), .B(n202), .ZN(n9) );
  OAOI211V2_8TH40 U7 ( .A1(n154), .A2(n136), .B(n153), .C(n196), .ZN(n14) );
  OAI211V2_8TH40 U8 ( .A1(n39), .A2(n17), .B(n197), .C(n208), .ZN(n45) );
  OAI31V2_8TH40 U9 ( .A1(n276), .A2(n40), .A3(n206), .B(n1), .ZN(n271) );
  OAI31V2_8TH40 U10 ( .A1(n350), .A2(n204), .A3(n206), .B(n277), .ZN(n217) );
  I2NOR4V2_8TH40 U11 ( .A1(n115), .A2(n263), .B1(n153), .B2(n40), .ZN(n254) );
  OAI22V2_8TH40 U12 ( .A1(n215), .A2(n216), .B1(n210), .B2(n218), .ZN(
        except_type_o[0]) );
  AOI31V2_8TH40 U13 ( .A1(n315), .A2(n268), .A3(n262), .B(rst), .ZN(n305) );
  OAI21V2_8TH40 U14 ( .A1(n236), .A2(n237), .B(n352), .ZN(n215) );
  NAND4V2_8TH40 U15 ( .A1(n242), .A2(n243), .A3(n244), .A4(n245), .ZN(n236) );
  NAND4V2_8TH40 U16 ( .A1(n238), .A2(n239), .A3(n240), .A4(n241), .ZN(n237) );
  OAI211V2_8TH40 U17 ( .A1(n6), .A2(n20), .B(n21), .C(n22), .ZN(
        exe_result_o[8]) );
  AOI21V2_8TH40 U18 ( .A1(n1), .A2(n23), .B(n13), .ZN(n21) );
  OAI211V2_8TH40 U19 ( .A1(n6), .A2(n185), .B(n186), .C(n187), .ZN(
        exe_result_o[10]) );
  AOI21V2_8TH40 U20 ( .A1(n1), .A2(n190), .B(n13), .ZN(n186) );
  OAI211V2_8TH40 U21 ( .A1(n6), .A2(n180), .B(n181), .C(n182), .ZN(
        exe_result_o[11]) );
  AOI21V2_8TH40 U22 ( .A1(n1), .A2(n183), .B(n13), .ZN(n181) );
  OAI211V2_8TH40 U23 ( .A1(n6), .A2(n175), .B(n176), .C(n177), .ZN(
        exe_result_o[12]) );
  AOI21V2_8TH40 U24 ( .A1(n1), .A2(n178), .B(n13), .ZN(n176) );
  OAI211V2_8TH40 U25 ( .A1(n6), .A2(n170), .B(n171), .C(n172), .ZN(
        exe_result_o[13]) );
  AOI21V2_8TH40 U26 ( .A1(n1), .A2(n173), .B(n13), .ZN(n171) );
  OAI211V2_8TH40 U27 ( .A1(n6), .A2(n165), .B(n166), .C(n167), .ZN(
        exe_result_o[14]) );
  AOI21V2_8TH40 U28 ( .A1(n1), .A2(n168), .B(n13), .ZN(n166) );
  OAI211V2_8TH40 U29 ( .A1(n5), .A2(n6), .B(n7), .C(n8), .ZN(exe_result_o[9])
         );
  AOI21V2_8TH40 U30 ( .A1(n1), .A2(n12), .B(n13), .ZN(n7) );
  OAI211V2_8TH40 U31 ( .A1(n155), .A2(n6), .B(n156), .C(n157), .ZN(
        exe_result_o[15]) );
  AOI21V2_8TH40 U32 ( .A1(n1), .A2(n158), .B(n69), .ZN(n156) );
  OAI211V2_8TH40 U33 ( .A1(n60), .A2(n4), .B(n61), .C(n62), .ZN(
        exe_result_o[31]) );
  OAI211V2_8TH40 U34 ( .A1(n220), .A2(n221), .B(n222), .C(n223), .ZN(n216) );
  OAI211V2_8TH40 U35 ( .A1(n26), .A2(n65), .B(n109), .C(n110), .ZN(
        exe_result_o[24]) );
  AOI21V2_8TH40 U36 ( .A1(n1), .A2(n111), .B(n69), .ZN(n109) );
  OAI211V2_8TH40 U37 ( .A1(n16), .A2(n65), .B(n104), .C(n105), .ZN(
        exe_result_o[25]) );
  AOI21V2_8TH40 U38 ( .A1(n1), .A2(n106), .B(n69), .ZN(n104) );
  OAI211V2_8TH40 U39 ( .A1(n79), .A2(n65), .B(n98), .C(n99), .ZN(
        exe_result_o[26]) );
  AOI21V2_8TH40 U40 ( .A1(n1), .A2(n100), .B(n69), .ZN(n98) );
  OAI211V2_8TH40 U41 ( .A1(n59), .A2(n65), .B(n92), .C(n93), .ZN(
        exe_result_o[27]) );
  AOI21V2_8TH40 U42 ( .A1(n1), .A2(n94), .B(n69), .ZN(n92) );
  OAI211V2_8TH40 U43 ( .A1(n55), .A2(n65), .B(n86), .C(n87), .ZN(
        exe_result_o[28]) );
  AOI21V2_8TH40 U44 ( .A1(n1), .A2(n88), .B(n69), .ZN(n86) );
  OAI211V2_8TH40 U45 ( .A1(n51), .A2(n65), .B(n80), .C(n81), .ZN(
        exe_result_o[29]) );
  AOI21V2_8TH40 U46 ( .A1(n1), .A2(n82), .B(n69), .ZN(n80) );
  OAI211V2_8TH40 U47 ( .A1(n47), .A2(n65), .B(n66), .C(n67), .ZN(
        exe_result_o[30]) );
  AOI21V2_8TH40 U48 ( .A1(n1), .A2(n68), .B(n69), .ZN(n66) );
  AOAI211V2_8TH40 U49 ( .A1(n48), .A2(n49), .B(n4), .C(n50), .ZN(
        exe_result_o[5]) );
  AOAI211V2_8TH40 U50 ( .A1(n41), .A2(n42), .B(n4), .C(n43), .ZN(
        exe_result_o[6]) );
  AOAI211V2_8TH40 U51 ( .A1(n198), .A2(n199), .B(n4), .C(n200), .ZN(
        exe_result_o[0]) );
  AOAI211V2_8TH40 U52 ( .A1(n133), .A2(n134), .B(n4), .C(n135), .ZN(
        exe_result_o[1]) );
  AOAI211V2_8TH40 U53 ( .A1(n76), .A2(n77), .B(n4), .C(n78), .ZN(
        exe_result_o[2]) );
  AOAI211V2_8TH40 U54 ( .A1(n56), .A2(n57), .B(n4), .C(n58), .ZN(
        exe_result_o[3]) );
  AOAI211V2_8TH40 U55 ( .A1(n52), .A2(n53), .B(n4), .C(n54), .ZN(
        exe_result_o[4]) );
  OAI222V2_8TH40 U56 ( .A1(n161), .A2(n17), .B1(n14), .B2(n163), .C1(n164), 
        .C2(n19), .ZN(n158) );
  OAI221V2_8TH40 U57 ( .A1(n25), .A2(n250), .B1(n113), .B2(n303), .C(n313), 
        .ZN(N586) );
  OAI221V2_8TH40 U58 ( .A1(n15), .A2(n250), .B1(n108), .B2(n303), .C(n312), 
        .ZN(N587) );
  OAI221V2_8TH40 U59 ( .A1(n193), .A2(n250), .B1(n102), .B2(n303), .C(n311), 
        .ZN(N588) );
  OAI221V2_8TH40 U60 ( .A1(n184), .A2(n250), .B1(n96), .B2(n303), .C(n310), 
        .ZN(N589) );
  OAI221V2_8TH40 U61 ( .A1(n179), .A2(n250), .B1(n90), .B2(n303), .C(n309), 
        .ZN(N590) );
  OAI221V2_8TH40 U62 ( .A1(n174), .A2(n250), .B1(n84), .B2(n303), .C(n308), 
        .ZN(N591) );
  OAI221V2_8TH40 U63 ( .A1(n169), .A2(n250), .B1(n73), .B2(n303), .C(n307), 
        .ZN(N592) );
  OAI221V2_8TH40 U64 ( .A1(n163), .A2(n250), .B1(n283), .B2(n303), .C(n304), 
        .ZN(N593) );
  OAI221V2_8TH40 U65 ( .A1(n25), .A2(n303), .B1(n301), .B2(n337), .C(n347), 
        .ZN(N570) );
  OAI221V2_8TH40 U66 ( .A1(n15), .A2(n303), .B1(n299), .B2(n337), .C(n346), 
        .ZN(N571) );
  OAI221V2_8TH40 U67 ( .A1(n193), .A2(n303), .B1(n297), .B2(n337), .C(n345), 
        .ZN(N572) );
  OAI221V2_8TH40 U68 ( .A1(n184), .A2(n303), .B1(n295), .B2(n337), .C(n344), 
        .ZN(N573) );
  OAI221V2_8TH40 U69 ( .A1(n179), .A2(n303), .B1(n293), .B2(n337), .C(n343), 
        .ZN(N574) );
  OAI221V2_8TH40 U70 ( .A1(n174), .A2(n303), .B1(n291), .B2(n337), .C(n342), 
        .ZN(N575) );
  OAI221V2_8TH40 U71 ( .A1(n169), .A2(n303), .B1(n289), .B2(n337), .C(n341), 
        .ZN(N576) );
  OAI221V2_8TH40 U72 ( .A1(n163), .A2(n303), .B1(n285), .B2(n337), .C(n338), 
        .ZN(N577) );
  OAI221V2_8TH40 U73 ( .A1(n113), .A2(n284), .B1(n301), .B2(n250), .C(n302), 
        .ZN(N594) );
  OAI221V2_8TH40 U74 ( .A1(n108), .A2(n284), .B1(n299), .B2(n250), .C(n300), 
        .ZN(N595) );
  OAI221V2_8TH40 U75 ( .A1(n102), .A2(n284), .B1(n297), .B2(n250), .C(n298), 
        .ZN(N596) );
  OAI221V2_8TH40 U76 ( .A1(n96), .A2(n284), .B1(n295), .B2(n250), .C(n296), 
        .ZN(N597) );
  OAI221V2_8TH40 U77 ( .A1(n90), .A2(n284), .B1(n293), .B2(n250), .C(n294), 
        .ZN(N598) );
  OAI221V2_8TH40 U78 ( .A1(n84), .A2(n284), .B1(n291), .B2(n250), .C(n292), 
        .ZN(N599) );
  OAI221V2_8TH40 U79 ( .A1(n73), .A2(n284), .B1(n289), .B2(n250), .C(n290), 
        .ZN(N600) );
  OAI221V2_8TH40 U80 ( .A1(n283), .A2(n284), .B1(n285), .B2(n250), .C(n286), 
        .ZN(N601) );
  OAI22V2_8TH40 U81 ( .A1(n191), .A2(n265), .B1(n266), .B2(n267), .ZN(n205) );
  OAI221V2_8TH40 U82 ( .A1(n316), .A2(n335), .B1(n25), .B2(n318), .C(n336), 
        .ZN(N578) );
  OAI221V2_8TH40 U83 ( .A1(n316), .A2(n332), .B1(n15), .B2(n318), .C(n334), 
        .ZN(N579) );
  OAI221V2_8TH40 U84 ( .A1(n316), .A2(n330), .B1(n193), .B2(n318), .C(n331), 
        .ZN(N580) );
  OAI221V2_8TH40 U85 ( .A1(n316), .A2(n328), .B1(n184), .B2(n318), .C(n329), 
        .ZN(N581) );
  OAI221V2_8TH40 U86 ( .A1(n316), .A2(n326), .B1(n179), .B2(n318), .C(n327), 
        .ZN(N582) );
  OAI221V2_8TH40 U87 ( .A1(n316), .A2(n324), .B1(n174), .B2(n318), .C(n325), 
        .ZN(N583) );
  OAI221V2_8TH40 U88 ( .A1(n316), .A2(n322), .B1(n169), .B2(n318), .C(n323), 
        .ZN(N584) );
  OAI221V2_8TH40 U89 ( .A1(n316), .A2(n317), .B1(n163), .B2(n318), .C(n319), 
        .ZN(N585) );
  OAI21V2_8TH40 U90 ( .A1(n159), .A2(n160), .B(n1), .ZN(n61) );
  AOI211V2_8TH40 U91 ( .A1(wb_cp0_wdata[15]), .A2(cp0_cause[15]), .B(n227), 
        .C(n228), .ZN(n226) );
  AOI21V2_8TH40 U92 ( .A1(n203), .A2(n256), .B(n257), .ZN(n251) );
  NAND2V2_8TH40 U93 ( .A1(n145), .A2(n146), .ZN(exe_result_o[17]) );
  AOI211V2_8TH40 U94 ( .A1(ls_data_tmp[17]), .A2(n118), .B(n147), .C(n69), 
        .ZN(n146) );
  OAI22V2_8TH40 U95 ( .A1(n6), .A2(n148), .B1(n107), .B2(n120), .ZN(n147) );
  NAND2V2_8TH40 U96 ( .A1(n116), .A2(n117), .ZN(exe_result_o[23]) );
  AOI211V2_8TH40 U97 ( .A1(ls_data_tmp[23]), .A2(n118), .B(n119), .C(n69), 
        .ZN(n117) );
  OAI211V2_8TH40 U98 ( .A1(rst), .A2(n249), .B(n250), .C(n251), .ZN(
        dmem_byte_sel[2]) );
  AOAI211V2_8TH40 U99 ( .A1(n246), .A2(n247), .B(rst), .C(n202), .ZN(
        dmem_byte_sel[3]) );
  NAND2V2_8TH40 U100 ( .A1(n213), .A2(n214), .ZN(except_type_o[1]) );
  IOA21V2_8TH40 U101 ( .A1(exe_result[7]), .A2(n9), .B(n27), .ZN(
        exe_result_o[7]) );
  AOI32V2_8TH40 U102 ( .A1(dmem_data_i[7]), .A2(n28), .A3(n29), .B1(n1), .B2(
        n30), .ZN(n27) );
  AO221V2_8TH40 U103 ( .A1(n31), .A2(n32), .B1(n33), .B2(ls_data_tmp[7]), .C(
        n34), .Z(n30) );
  OAI32V2_8TH40 U104 ( .A1(n35), .A2(n36), .A3(n17), .B1(n37), .B2(n38), .ZN(
        n34) );
  NAND2V2_8TH40 U105 ( .A1(n149), .A2(n150), .ZN(exe_result_o[16]) );
  AOI211V2_8TH40 U106 ( .A1(ls_data_tmp[16]), .A2(n118), .B(n151), .C(n69), 
        .ZN(n150) );
  OAI22V2_8TH40 U107 ( .A1(n6), .A2(n152), .B1(n112), .B2(n120), .ZN(n151) );
  NAND2V2_8TH40 U108 ( .A1(n141), .A2(n142), .ZN(exe_result_o[18]) );
  AOI211V2_8TH40 U109 ( .A1(ls_data_tmp[18]), .A2(n118), .B(n143), .C(n69), 
        .ZN(n142) );
  OAI22V2_8TH40 U110 ( .A1(n6), .A2(n144), .B1(n101), .B2(n120), .ZN(n143) );
  NAND2V2_8TH40 U111 ( .A1(n137), .A2(n138), .ZN(exe_result_o[19]) );
  AOI211V2_8TH40 U112 ( .A1(ls_data_tmp[19]), .A2(n118), .B(n139), .C(n69), 
        .ZN(n138) );
  OAI22V2_8TH40 U113 ( .A1(n6), .A2(n140), .B1(n95), .B2(n120), .ZN(n139) );
  NAND2V2_8TH40 U114 ( .A1(n129), .A2(n130), .ZN(exe_result_o[20]) );
  AOI211V2_8TH40 U115 ( .A1(ls_data_tmp[20]), .A2(n118), .B(n131), .C(n69), 
        .ZN(n130) );
  OAI22V2_8TH40 U116 ( .A1(n6), .A2(n132), .B1(n89), .B2(n120), .ZN(n131) );
  NAND2V2_8TH40 U117 ( .A1(n125), .A2(n126), .ZN(exe_result_o[21]) );
  AOI211V2_8TH40 U118 ( .A1(ls_data_tmp[21]), .A2(n118), .B(n127), .C(n69), 
        .ZN(n126) );
  OAI22V2_8TH40 U119 ( .A1(n6), .A2(n128), .B1(n83), .B2(n120), .ZN(n127) );
  NAND2V2_8TH40 U120 ( .A1(n121), .A2(n122), .ZN(exe_result_o[22]) );
  AOI211V2_8TH40 U121 ( .A1(ls_data_tmp[22]), .A2(n118), .B(n123), .C(n69), 
        .ZN(n122) );
  OAI22V2_8TH40 U122 ( .A1(n6), .A2(n124), .B1(n70), .B2(n120), .ZN(n123) );
  INAND2V2_8TH40 U123 ( .A1(n348), .B1(n351), .ZN(n207) );
  INOR2V0_8TH40 U124 ( .A1(target_gpr[4]), .B1(rst), .ZN(target_gpr_o[4]) );
  INOR2V0_8TH40 U125 ( .A1(target_gpr[3]), .B1(rst), .ZN(target_gpr_o[3]) );
  INOR2V0_8TH40 U126 ( .A1(target_gpr[2]), .B1(rst), .ZN(target_gpr_o[2]) );
  INOR2V0_8TH40 U127 ( .A1(target_gpr[1]), .B1(rst), .ZN(target_gpr_o[1]) );
  INOR2V0_8TH40 U128 ( .A1(target_gpr[0]), .B1(rst), .ZN(target_gpr_o[0]) );
  AO21V0_8TH40 U129 ( .A1(n1), .A2(n2), .B(mem_llbit_value), .Z(mem_llbit_we)
         );
  NOR2V0P5_8TH40 U130 ( .A1(n3), .A2(n4), .ZN(mem_llbit_value) );
  INOR2V0_8TH40 U131 ( .A1(lo[9]), .B1(rst), .ZN(lo_o[9]) );
  INOR2V0_8TH40 U132 ( .A1(lo[8]), .B1(rst), .ZN(lo_o[8]) );
  INOR2V0_8TH40 U133 ( .A1(lo[7]), .B1(rst), .ZN(lo_o[7]) );
  INOR2V0_8TH40 U134 ( .A1(lo[6]), .B1(rst), .ZN(lo_o[6]) );
  INOR2V0_8TH40 U135 ( .A1(lo[5]), .B1(rst), .ZN(lo_o[5]) );
  INOR2V0_8TH40 U136 ( .A1(lo[4]), .B1(rst), .ZN(lo_o[4]) );
  INOR2V0_8TH40 U137 ( .A1(lo[3]), .B1(rst), .ZN(lo_o[3]) );
  INOR2V0_8TH40 U138 ( .A1(lo[31]), .B1(rst), .ZN(lo_o[31]) );
  INOR2V0_8TH40 U139 ( .A1(lo[30]), .B1(rst), .ZN(lo_o[30]) );
  INOR2V0_8TH40 U140 ( .A1(lo[2]), .B1(rst), .ZN(lo_o[2]) );
  INOR2V0_8TH40 U141 ( .A1(lo[29]), .B1(rst), .ZN(lo_o[29]) );
  INOR2V0_8TH40 U142 ( .A1(lo[28]), .B1(rst), .ZN(lo_o[28]) );
  INOR2V0_8TH40 U143 ( .A1(lo[27]), .B1(rst), .ZN(lo_o[27]) );
  INOR2V0_8TH40 U144 ( .A1(lo[26]), .B1(rst), .ZN(lo_o[26]) );
  INOR2V0_8TH40 U145 ( .A1(lo[25]), .B1(rst), .ZN(lo_o[25]) );
  INOR2V0_8TH40 U146 ( .A1(lo[24]), .B1(rst), .ZN(lo_o[24]) );
  INOR2V0_8TH40 U147 ( .A1(lo[23]), .B1(rst), .ZN(lo_o[23]) );
  INOR2V0_8TH40 U148 ( .A1(lo[22]), .B1(rst), .ZN(lo_o[22]) );
  INOR2V0_8TH40 U149 ( .A1(lo[21]), .B1(rst), .ZN(lo_o[21]) );
  INOR2V0_8TH40 U150 ( .A1(lo[20]), .B1(rst), .ZN(lo_o[20]) );
  INOR2V0_8TH40 U151 ( .A1(lo[1]), .B1(rst), .ZN(lo_o[1]) );
  INOR2V0_8TH40 U152 ( .A1(lo[19]), .B1(rst), .ZN(lo_o[19]) );
  INOR2V0_8TH40 U153 ( .A1(lo[18]), .B1(rst), .ZN(lo_o[18]) );
  INOR2V0_8TH40 U154 ( .A1(lo[17]), .B1(rst), .ZN(lo_o[17]) );
  INOR2V0_8TH40 U155 ( .A1(lo[16]), .B1(rst), .ZN(lo_o[16]) );
  INOR2V0_8TH40 U156 ( .A1(lo[15]), .B1(rst), .ZN(lo_o[15]) );
  INOR2V0_8TH40 U157 ( .A1(lo[14]), .B1(rst), .ZN(lo_o[14]) );
  INOR2V0_8TH40 U158 ( .A1(lo[13]), .B1(rst), .ZN(lo_o[13]) );
  INOR2V0_8TH40 U159 ( .A1(lo[12]), .B1(rst), .ZN(lo_o[12]) );
  INOR2V0_8TH40 U160 ( .A1(lo[11]), .B1(rst), .ZN(lo_o[11]) );
  INOR2V0_8TH40 U161 ( .A1(lo[10]), .B1(rst), .ZN(lo_o[10]) );
  INOR2V0_8TH40 U162 ( .A1(lo[0]), .B1(rst), .ZN(lo_o[0]) );
  INOR2V0_8TH40 U163 ( .A1(hilo_we), .B1(rst), .ZN(hilo_we_o) );
  INOR2V0_8TH40 U164 ( .A1(hi[9]), .B1(rst), .ZN(hi_o[9]) );
  INOR2V0_8TH40 U165 ( .A1(hi[8]), .B1(rst), .ZN(hi_o[8]) );
  INOR2V0_8TH40 U166 ( .A1(hi[7]), .B1(rst), .ZN(hi_o[7]) );
  INOR2V0_8TH40 U167 ( .A1(hi[6]), .B1(rst), .ZN(hi_o[6]) );
  INOR2V0_8TH40 U168 ( .A1(hi[5]), .B1(rst), .ZN(hi_o[5]) );
  INOR2V0_8TH40 U169 ( .A1(hi[4]), .B1(rst), .ZN(hi_o[4]) );
  INOR2V0_8TH40 U170 ( .A1(hi[3]), .B1(rst), .ZN(hi_o[3]) );
  INOR2V0_8TH40 U171 ( .A1(hi[31]), .B1(rst), .ZN(hi_o[31]) );
  INOR2V0_8TH40 U172 ( .A1(hi[30]), .B1(rst), .ZN(hi_o[30]) );
  INOR2V0_8TH40 U173 ( .A1(hi[2]), .B1(rst), .ZN(hi_o[2]) );
  INOR2V0_8TH40 U174 ( .A1(hi[29]), .B1(rst), .ZN(hi_o[29]) );
  INOR2V0_8TH40 U175 ( .A1(hi[28]), .B1(rst), .ZN(hi_o[28]) );
  INOR2V0_8TH40 U176 ( .A1(hi[27]), .B1(rst), .ZN(hi_o[27]) );
  INOR2V0_8TH40 U177 ( .A1(hi[26]), .B1(rst), .ZN(hi_o[26]) );
  INOR2V0_8TH40 U178 ( .A1(hi[25]), .B1(rst), .ZN(hi_o[25]) );
  INOR2V0_8TH40 U179 ( .A1(hi[24]), .B1(rst), .ZN(hi_o[24]) );
  INOR2V0_8TH40 U180 ( .A1(hi[23]), .B1(rst), .ZN(hi_o[23]) );
  INOR2V0_8TH40 U181 ( .A1(hi[22]), .B1(rst), .ZN(hi_o[22]) );
  INOR2V0_8TH40 U182 ( .A1(hi[21]), .B1(rst), .ZN(hi_o[21]) );
  INOR2V0_8TH40 U183 ( .A1(hi[20]), .B1(rst), .ZN(hi_o[20]) );
  INOR2V0_8TH40 U184 ( .A1(hi[1]), .B1(rst), .ZN(hi_o[1]) );
  INOR2V0_8TH40 U185 ( .A1(hi[19]), .B1(rst), .ZN(hi_o[19]) );
  INOR2V0_8TH40 U186 ( .A1(hi[18]), .B1(rst), .ZN(hi_o[18]) );
  INOR2V0_8TH40 U187 ( .A1(hi[17]), .B1(rst), .ZN(hi_o[17]) );
  INOR2V0_8TH40 U188 ( .A1(hi[16]), .B1(rst), .ZN(hi_o[16]) );
  INOR2V0_8TH40 U189 ( .A1(hi[15]), .B1(rst), .ZN(hi_o[15]) );
  INOR2V0_8TH40 U190 ( .A1(hi[14]), .B1(rst), .ZN(hi_o[14]) );
  INOR2V0_8TH40 U191 ( .A1(hi[13]), .B1(rst), .ZN(hi_o[13]) );
  INOR2V0_8TH40 U192 ( .A1(hi[12]), .B1(rst), .ZN(hi_o[12]) );
  INOR2V0_8TH40 U193 ( .A1(hi[11]), .B1(rst), .ZN(hi_o[11]) );
  INOR2V0_8TH40 U194 ( .A1(hi[10]), .B1(rst), .ZN(hi_o[10]) );
  INOR2V0_8TH40 U195 ( .A1(hi[0]), .B1(rst), .ZN(hi_o[0]) );
  INOR2V0_8TH40 U196 ( .A1(gpr_we), .B1(rst), .ZN(gpr_we_o) );
  AOI222V0_8TH40 U197 ( .A1(exe_result[9]), .A2(n9), .B1(dmem_data_i[17]), 
        .B2(n10), .C1(dmem_data_i[1]), .C2(n11), .ZN(n8) );
  OAI222V0_8TH40 U198 ( .A1(n14), .A2(n15), .B1(n16), .B2(n17), .C1(n18), .C2(
        n19), .ZN(n12) );
  CLKNV1_8TH40 U199 ( .I(dmem_data_i[9]), .ZN(n5) );
  AOI222V0_8TH40 U200 ( .A1(exe_result[8]), .A2(n9), .B1(dmem_data_i[16]), 
        .B2(n10), .C1(dmem_data_i[0]), .C2(n11), .ZN(n22) );
  OAI222V0_8TH40 U201 ( .A1(n19), .A2(n24), .B1(n14), .B2(n25), .C1(n26), .C2(
        n17), .ZN(n23) );
  CLKNV1_8TH40 U202 ( .I(dmem_data_i[8]), .ZN(n20) );
  IAO21V0_8TH40 U203 ( .A1(n39), .A2(n17), .B(n40), .ZN(n38) );
  CLKNAND2V1_8TH40 U204 ( .A1(exe_result[6]), .A2(n9), .ZN(n43) );
  AOI22V0_8TH40 U205 ( .A1(dmem_data_i[22]), .A2(n44), .B1(dmem_data_i[6]), 
        .B2(n45), .ZN(n42) );
  IAO22V0_8TH40 U206 ( .B1(ls_data_tmp[6]), .B2(n33), .A1(n46), .A2(n47), .ZN(
        n41) );
  CLKNAND2V1_8TH40 U207 ( .A1(exe_result[5]), .A2(n9), .ZN(n50) );
  AOI22V0_8TH40 U208 ( .A1(dmem_data_i[21]), .A2(n44), .B1(dmem_data_i[5]), 
        .B2(n45), .ZN(n49) );
  IAO22V0_8TH40 U209 ( .B1(ls_data_tmp[5]), .B2(n33), .A1(n46), .A2(n51), .ZN(
        n48) );
  CLKNAND2V1_8TH40 U210 ( .A1(exe_result[4]), .A2(n9), .ZN(n54) );
  AOI22V0_8TH40 U211 ( .A1(dmem_data_i[20]), .A2(n44), .B1(dmem_data_i[4]), 
        .B2(n45), .ZN(n53) );
  IAO22V0_8TH40 U212 ( .B1(ls_data_tmp[4]), .B2(n33), .A1(n46), .A2(n55), .ZN(
        n52) );
  CLKNAND2V1_8TH40 U213 ( .A1(exe_result[3]), .A2(n9), .ZN(n58) );
  AOI22V0_8TH40 U214 ( .A1(dmem_data_i[19]), .A2(n44), .B1(dmem_data_i[3]), 
        .B2(n45), .ZN(n57) );
  IAO22V0_8TH40 U215 ( .B1(ls_data_tmp[3]), .B2(n33), .A1(n46), .A2(n59), .ZN(
        n56) );
  AOI22V0_8TH40 U216 ( .A1(n29), .A2(n31), .B1(exe_result[31]), .B2(n9), .ZN(
        n62) );
  AOI22V0_8TH40 U217 ( .A1(ls_data_tmp[31]), .A2(n63), .B1(dmem_data_i[31]), 
        .B2(n64), .ZN(n60) );
  AOI22V0_8TH40 U218 ( .A1(dmem_data_i[22]), .A2(n11), .B1(exe_result[30]), 
        .B2(n9), .ZN(n67) );
  OAI222V0_8TH40 U219 ( .A1(n70), .A2(n71), .B1(n72), .B2(n73), .C1(n74), .C2(
        n75), .ZN(n68) );
  CLKNAND2V1_8TH40 U220 ( .A1(exe_result[2]), .A2(n9), .ZN(n78) );
  AOI22V0_8TH40 U221 ( .A1(dmem_data_i[18]), .A2(n44), .B1(dmem_data_i[2]), 
        .B2(n45), .ZN(n77) );
  IAO22V0_8TH40 U222 ( .B1(ls_data_tmp[2]), .B2(n33), .A1(n46), .A2(n79), .ZN(
        n76) );
  AOI22V0_8TH40 U223 ( .A1(dmem_data_i[21]), .A2(n11), .B1(exe_result[29]), 
        .B2(n9), .ZN(n81) );
  OAI222V0_8TH40 U224 ( .A1(n83), .A2(n71), .B1(n72), .B2(n84), .C1(n74), .C2(
        n85), .ZN(n82) );
  AOI22V0_8TH40 U225 ( .A1(dmem_data_i[20]), .A2(n11), .B1(exe_result[28]), 
        .B2(n9), .ZN(n87) );
  OAI222V0_8TH40 U226 ( .A1(n89), .A2(n71), .B1(n72), .B2(n90), .C1(n74), .C2(
        n91), .ZN(n88) );
  AOI22V0_8TH40 U227 ( .A1(dmem_data_i[19]), .A2(n11), .B1(exe_result[27]), 
        .B2(n9), .ZN(n93) );
  OAI222V0_8TH40 U228 ( .A1(n95), .A2(n71), .B1(n72), .B2(n96), .C1(n74), .C2(
        n97), .ZN(n94) );
  AOI22V0_8TH40 U229 ( .A1(dmem_data_i[18]), .A2(n11), .B1(exe_result[26]), 
        .B2(n9), .ZN(n99) );
  OAI222V0_8TH40 U230 ( .A1(n71), .A2(n101), .B1(n72), .B2(n102), .C1(n74), 
        .C2(n103), .ZN(n100) );
  AOI22V0_8TH40 U231 ( .A1(n11), .A2(dmem_data_i[17]), .B1(exe_result[25]), 
        .B2(n9), .ZN(n105) );
  OAI222V0_8TH40 U232 ( .A1(n107), .A2(n71), .B1(n72), .B2(n108), .C1(n74), 
        .C2(n18), .ZN(n106) );
  CLKNV1_8TH40 U233 ( .I(dmem_data_i[25]), .ZN(n18) );
  AOI22V0_8TH40 U234 ( .A1(dmem_data_i[16]), .A2(n11), .B1(exe_result[24]), 
        .B2(n9), .ZN(n110) );
  OAI222V0_8TH40 U235 ( .A1(n112), .A2(n71), .B1(n72), .B2(n113), .C1(n74), 
        .C2(n24), .ZN(n111) );
  CLKNV1_8TH40 U236 ( .I(dmem_data_i[24]), .ZN(n24) );
  CLKNV1_8TH40 U237 ( .I(n64), .ZN(n74) );
  CLKNV1_8TH40 U238 ( .I(n63), .ZN(n72) );
  AOI21V0_8TH40 U239 ( .A1(n39), .A2(n114), .B(n115), .ZN(n63) );
  OAI22V0_8TH40 U240 ( .A1(n35), .A2(n6), .B1(n37), .B2(n120), .ZN(n119) );
  AOI222V0_8TH40 U241 ( .A1(exe_result[23]), .A2(n9), .B1(n10), .B2(
        dmem_data_i[31]), .C1(n11), .C2(dmem_data_i[15]), .ZN(n116) );
  CLKNV1_8TH40 U242 ( .I(dmem_data_i[6]), .ZN(n70) );
  CLKNV1_8TH40 U243 ( .I(dmem_data_i[22]), .ZN(n124) );
  AOI222V0_8TH40 U244 ( .A1(exe_result[22]), .A2(n9), .B1(dmem_data_i[30]), 
        .B2(n10), .C1(dmem_data_i[14]), .C2(n11), .ZN(n121) );
  CLKNV1_8TH40 U245 ( .I(dmem_data_i[5]), .ZN(n83) );
  CLKNV1_8TH40 U246 ( .I(dmem_data_i[21]), .ZN(n128) );
  AOI222V0_8TH40 U247 ( .A1(exe_result[21]), .A2(n9), .B1(dmem_data_i[29]), 
        .B2(n10), .C1(dmem_data_i[13]), .C2(n11), .ZN(n125) );
  CLKNV1_8TH40 U248 ( .I(dmem_data_i[4]), .ZN(n89) );
  CLKNV1_8TH40 U249 ( .I(dmem_data_i[20]), .ZN(n132) );
  AOI222V0_8TH40 U250 ( .A1(exe_result[20]), .A2(n9), .B1(dmem_data_i[28]), 
        .B2(n10), .C1(dmem_data_i[12]), .C2(n11), .ZN(n129) );
  CLKNAND2V1_8TH40 U251 ( .A1(exe_result[1]), .A2(n9), .ZN(n135) );
  AOI22V0_8TH40 U252 ( .A1(dmem_data_i[17]), .A2(n44), .B1(dmem_data_i[1]), 
        .B2(n45), .ZN(n134) );
  IAO22V0_8TH40 U253 ( .B1(ls_data_tmp[1]), .B2(n33), .A1(n46), .A2(n16), .ZN(
        n133) );
  AOI22V0_8TH40 U254 ( .A1(n136), .A2(dmem_data_i[9]), .B1(n28), .B2(
        dmem_data_i[25]), .ZN(n16) );
  CLKNV1_8TH40 U255 ( .I(dmem_data_i[3]), .ZN(n95) );
  CLKNV1_8TH40 U256 ( .I(dmem_data_i[19]), .ZN(n140) );
  AOI222V0_8TH40 U257 ( .A1(exe_result[19]), .A2(n9), .B1(dmem_data_i[27]), 
        .B2(n10), .C1(dmem_data_i[11]), .C2(n11), .ZN(n137) );
  CLKNV1_8TH40 U258 ( .I(dmem_data_i[2]), .ZN(n101) );
  CLKNV1_8TH40 U259 ( .I(dmem_data_i[18]), .ZN(n144) );
  AOI222V0_8TH40 U260 ( .A1(exe_result[18]), .A2(n9), .B1(dmem_data_i[26]), 
        .B2(n10), .C1(dmem_data_i[10]), .C2(n11), .ZN(n141) );
  CLKNV1_8TH40 U261 ( .I(dmem_data_i[1]), .ZN(n107) );
  CLKNV1_8TH40 U262 ( .I(dmem_data_i[17]), .ZN(n148) );
  AOI222V0_8TH40 U263 ( .A1(exe_result[17]), .A2(n9), .B1(n10), .B2(
        dmem_data_i[25]), .C1(n11), .C2(dmem_data_i[9]), .ZN(n145) );
  CLKNAND2V1_8TH40 U264 ( .A1(n29), .A2(n136), .ZN(n120) );
  CLKNV1_8TH40 U265 ( .I(n65), .ZN(n29) );
  CLKNV1_8TH40 U266 ( .I(dmem_data_i[0]), .ZN(n112) );
  CLKNV1_8TH40 U267 ( .I(dmem_data_i[16]), .ZN(n152) );
  OAOI211V0_8TH40 U268 ( .A1(n115), .A2(n114), .B(n71), .C(n4), .ZN(n118) );
  CLKNAND2V1_8TH40 U269 ( .A1(n153), .A2(n154), .ZN(n71) );
  AOI222V0_8TH40 U270 ( .A1(exe_result[16]), .A2(n9), .B1(dmem_data_i[24]), 
        .B2(n10), .C1(dmem_data_i[8]), .C2(n11), .ZN(n149) );
  AOI222V0_8TH40 U271 ( .A1(exe_result[15]), .A2(n9), .B1(n10), .B2(
        dmem_data_i[23]), .C1(n11), .C2(dmem_data_i[7]), .ZN(n157) );
  CLKNV1_8TH40 U272 ( .I(n61), .ZN(n69) );
  NOR4V0P5_8TH40 U273 ( .A1(inst_type[3]), .A2(inst_type[1]), .A3(n161), .A4(
        n162), .ZN(n159) );
  CLKNV1_8TH40 U274 ( .I(dmem_data_i[31]), .ZN(n164) );
  CLKNV1_8TH40 U275 ( .I(dmem_data_i[15]), .ZN(n155) );
  AOI222V0_8TH40 U276 ( .A1(exe_result[14]), .A2(n9), .B1(dmem_data_i[22]), 
        .B2(n10), .C1(dmem_data_i[6]), .C2(n11), .ZN(n167) );
  OAI222V0_8TH40 U277 ( .A1(n14), .A2(n169), .B1(n47), .B2(n17), .C1(n19), 
        .C2(n75), .ZN(n168) );
  CLKNV1_8TH40 U278 ( .I(dmem_data_i[30]), .ZN(n75) );
  AOI22V0_8TH40 U279 ( .A1(n28), .A2(dmem_data_i[30]), .B1(n136), .B2(
        dmem_data_i[14]), .ZN(n47) );
  CLKNV1_8TH40 U280 ( .I(dmem_data_i[14]), .ZN(n165) );
  AOI222V0_8TH40 U281 ( .A1(exe_result[13]), .A2(n9), .B1(dmem_data_i[21]), 
        .B2(n10), .C1(dmem_data_i[5]), .C2(n11), .ZN(n172) );
  OAI222V0_8TH40 U282 ( .A1(n14), .A2(n174), .B1(n51), .B2(n17), .C1(n19), 
        .C2(n85), .ZN(n173) );
  CLKNV1_8TH40 U283 ( .I(dmem_data_i[29]), .ZN(n85) );
  AOI22V0_8TH40 U284 ( .A1(n28), .A2(dmem_data_i[29]), .B1(n136), .B2(
        dmem_data_i[13]), .ZN(n51) );
  CLKNV1_8TH40 U285 ( .I(dmem_data_i[13]), .ZN(n170) );
  AOI222V0_8TH40 U286 ( .A1(exe_result[12]), .A2(n9), .B1(dmem_data_i[20]), 
        .B2(n10), .C1(dmem_data_i[4]), .C2(n11), .ZN(n177) );
  OAI222V0_8TH40 U287 ( .A1(n14), .A2(n179), .B1(n55), .B2(n17), .C1(n19), 
        .C2(n91), .ZN(n178) );
  CLKNV1_8TH40 U288 ( .I(dmem_data_i[28]), .ZN(n91) );
  AOI22V0_8TH40 U289 ( .A1(n28), .A2(dmem_data_i[28]), .B1(n136), .B2(
        dmem_data_i[12]), .ZN(n55) );
  CLKNV1_8TH40 U290 ( .I(dmem_data_i[12]), .ZN(n175) );
  AOI222V0_8TH40 U291 ( .A1(exe_result[11]), .A2(n9), .B1(dmem_data_i[19]), 
        .B2(n10), .C1(dmem_data_i[3]), .C2(n11), .ZN(n182) );
  OAI222V0_8TH40 U292 ( .A1(n14), .A2(n184), .B1(n59), .B2(n17), .C1(n19), 
        .C2(n97), .ZN(n183) );
  CLKNV1_8TH40 U293 ( .I(dmem_data_i[27]), .ZN(n97) );
  AOI22V0_8TH40 U294 ( .A1(n28), .A2(dmem_data_i[27]), .B1(n136), .B2(
        dmem_data_i[11]), .ZN(n59) );
  CLKNV1_8TH40 U295 ( .I(dmem_data_i[11]), .ZN(n180) );
  AOI222V0_8TH40 U296 ( .A1(exe_result[10]), .A2(n9), .B1(dmem_data_i[18]), 
        .B2(n10), .C1(dmem_data_i[2]), .C2(n11), .ZN(n187) );
  NOR3V0P5_8TH40 U297 ( .A1(n188), .A2(n4), .A3(n189), .ZN(n11) );
  NOR3V0P5_8TH40 U298 ( .A1(n39), .A2(n4), .A3(n115), .ZN(n10) );
  INOR2V0_8TH40 U299 ( .A1(n160), .B1(n4), .ZN(n13) );
  I2NOR4V0_8TH40 U300 ( .A1(n191), .A2(n31), .B1(inst_type[3]), .B2(
        inst_type[4]), .ZN(n160) );
  OAI221V0_8TH40 U301 ( .A1(n192), .A2(n37), .B1(n188), .B2(n35), .C(n161), 
        .ZN(n31) );
  AOI22V0_8TH40 U302 ( .A1(n28), .A2(dmem_data_i[31]), .B1(n136), .B2(
        dmem_data_i[15]), .ZN(n161) );
  CLKNV1_8TH40 U303 ( .I(dmem_data_i[23]), .ZN(n35) );
  CLKNV1_8TH40 U304 ( .I(dmem_data_i[7]), .ZN(n37) );
  OAI222V0_8TH40 U305 ( .A1(n14), .A2(n193), .B1(n79), .B2(n17), .C1(n19), 
        .C2(n103), .ZN(n190) );
  CLKNV1_8TH40 U306 ( .I(dmem_data_i[26]), .ZN(n103) );
  CLKNAND2V1_8TH40 U307 ( .A1(n194), .A2(n195), .ZN(n19) );
  AOI22V0_8TH40 U308 ( .A1(n28), .A2(dmem_data_i[26]), .B1(n136), .B2(
        dmem_data_i[10]), .ZN(n79) );
  NOR2V0P5_8TH40 U309 ( .A1(n115), .A2(n36), .ZN(n196) );
  CLKNV1_8TH40 U310 ( .I(dmem_data_i[10]), .ZN(n185) );
  AOAI211V0_8TH40 U311 ( .A1(n153), .A2(n28), .B(n64), .C(n1), .ZN(n6) );
  OAI21V0_8TH40 U312 ( .A1(n192), .A2(n115), .B(n197), .ZN(n64) );
  CLKNAND2V1_8TH40 U313 ( .A1(exe_result[0]), .A2(n9), .ZN(n200) );
  NOR4V0P5_8TH40 U314 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(n201)
         );
  AOI221V0_8TH40 U315 ( .A1(dmem_data_i[0]), .A2(n45), .B1(dmem_data_i[16]), 
        .B2(n44), .C(n2), .ZN(n199) );
  CLKNV1_8TH40 U316 ( .I(n207), .ZN(n2) );
  OAI22V0_8TH40 U317 ( .A1(n36), .A2(n17), .B1(n46), .B2(n188), .ZN(n44) );
  AOI22V0_8TH40 U318 ( .A1(n154), .A2(n32), .B1(n153), .B2(n28), .ZN(n208) );
  CLKNV1_8TH40 U319 ( .I(n192), .ZN(n154) );
  CLKNV1_8TH40 U320 ( .I(n40), .ZN(n197) );
  IAO22V0_8TH40 U321 ( .B1(ls_data_tmp[0]), .B2(n33), .A1(n46), .A2(n26), .ZN(
        n198) );
  AOI22V0_8TH40 U322 ( .A1(n136), .A2(dmem_data_i[8]), .B1(n28), .B2(
        dmem_data_i[24]), .ZN(n26) );
  CLKNV1_8TH40 U323 ( .I(n32), .ZN(n46) );
  CLKNAND2V1_8TH40 U324 ( .A1(n209), .A2(n115), .ZN(n32) );
  AOI31V0_8TH40 U325 ( .A1(n192), .A2(n188), .A3(n39), .B(n189), .ZN(n33) );
  OAI31V0_8TH40 U326 ( .A1(n210), .A2(n211), .A3(n212), .B(n213), .ZN(
        except_type_o[2]) );
  I2NAND4V0_8TH40 U327 ( .A1(except_type_i[8]), .A2(n215), .B1(
        except_type_i[9]), .B2(n216), .ZN(n214) );
  NOR4V0P5_8TH40 U328 ( .A1(rst), .A2(except_type_o[3]), .A3(except_type_o[0]), 
        .A4(n217), .ZN(dmem_we) );
  CLKNV1_8TH40 U329 ( .I(except_type_i[10]), .ZN(n218) );
  OR3V0_8TH40 U330 ( .A1(except_type_i[9]), .A2(except_type_i[8]), .A3(n215), 
        .Z(n210) );
  OAI31V0_8TH40 U331 ( .A1(n215), .A2(n211), .A3(n219), .B(n213), .ZN(
        except_type_o[3]) );
  I2NAND4V0_8TH40 U332 ( .A1(n215), .A2(n211), .B1(except_type_i[12]), .B2(
        n219), .ZN(n213) );
  INOR3V0_8TH40 U333 ( .A1(n212), .B1(except_type_i[8]), .B2(except_type_i[9]), 
        .ZN(n219) );
  NOR2V0P5_8TH40 U334 ( .A1(except_type_i[11]), .A2(except_type_i[10]), .ZN(
        n212) );
  CLKNV1_8TH40 U335 ( .I(n216), .ZN(n211) );
  MUX2NV0_8TH40 U336 ( .I0(cp0_status_i[1]), .I1(wb_cp0_wdata[1]), .S(n224), 
        .ZN(n223) );
  CKMUX2V2_8TH40 U337 ( .I0(cp0_status_i[0]), .I1(wb_cp0_wdata[0]), .S(n224), 
        .Z(n222) );
  MUX2NV0_8TH40 U338 ( .I0(n225), .I1(n226), .S(n224), .ZN(n221) );
  AO22V0_8TH40 U339 ( .A1(cp0_cause[14]), .A2(wb_cp0_wdata[14]), .B1(
        cp0_cause[13]), .B2(wb_cp0_wdata[13]), .Z(n228) );
  AO222V0_8TH40 U340 ( .A1(cp0_cause[11]), .A2(wb_cp0_wdata[11]), .B1(
        cp0_cause[10]), .B2(wb_cp0_wdata[10]), .C1(cp0_cause[12]), .C2(
        wb_cp0_wdata[12]), .Z(n227) );
  AOI222V0_8TH40 U341 ( .A1(cp0_status_i[12]), .A2(cp0_cause[12]), .B1(
        cp0_status_i[10]), .B2(cp0_cause[10]), .C1(cp0_status_i[11]), .C2(
        cp0_cause[11]), .ZN(n230) );
  AOI222V0_8TH40 U342 ( .A1(cp0_status_i[15]), .A2(cp0_cause[15]), .B1(
        cp0_status_i[13]), .B2(cp0_cause[13]), .C1(cp0_status_i[14]), .C2(
        cp0_cause[14]), .ZN(n229) );
  MUX2NV0_8TH40 U343 ( .I0(n231), .I1(n232), .S(n333), .ZN(n220) );
  I2NAND3V1_8TH40 U344 ( .A1(wb_cp0_waddr[1]), .A2(n233), .B(wb_cp0_waddr[0]), 
        .ZN(n333) );
  AOI22V0_8TH40 U345 ( .A1(cp0_cause_i[9]), .A2(n234), .B1(cp0_cause_i[8]), 
        .B2(n235), .ZN(n232) );
  AOI22V0_8TH40 U346 ( .A1(wb_cp0_wdata[9]), .A2(n234), .B1(wb_cp0_wdata[8]), 
        .B2(n235), .ZN(n231) );
  CKMUX2V2_8TH40 U347 ( .I0(cp0_status_i[8]), .I1(wb_cp0_wdata[8]), .S(n224), 
        .Z(n235) );
  CKMUX2V2_8TH40 U348 ( .I0(cp0_status_i[9]), .I1(wb_cp0_wdata[9]), .S(n224), 
        .Z(n234) );
  NOR3V0P5_8TH40 U349 ( .A1(wb_cp0_waddr[0]), .A2(wb_cp0_waddr[1]), .A3(n233), 
        .ZN(n224) );
  NOR4V0P5_8TH40 U350 ( .A1(cur_inst_addr_i[23]), .A2(cur_inst_addr_i[22]), 
        .A3(cur_inst_addr_i[21]), .A4(cur_inst_addr_i[20]), .ZN(n241) );
  NOR4V0P5_8TH40 U351 ( .A1(cur_inst_addr_i[1]), .A2(cur_inst_addr_i[19]), 
        .A3(cur_inst_addr_i[18]), .A4(cur_inst_addr_i[17]), .ZN(n240) );
  NOR4V0P5_8TH40 U352 ( .A1(cur_inst_addr_i[16]), .A2(cur_inst_addr_i[15]), 
        .A3(cur_inst_addr_i[14]), .A4(cur_inst_addr_i[13]), .ZN(n239) );
  NOR4V0P5_8TH40 U353 ( .A1(cur_inst_addr_i[12]), .A2(cur_inst_addr_i[11]), 
        .A3(cur_inst_addr_i[10]), .A4(cur_inst_addr_i[0]), .ZN(n238) );
  NOR4V0P5_8TH40 U354 ( .A1(cur_inst_addr_i[9]), .A2(cur_inst_addr_i[8]), .A3(
        cur_inst_addr_i[7]), .A4(cur_inst_addr_i[6]), .ZN(n245) );
  NOR4V0P5_8TH40 U355 ( .A1(cur_inst_addr_i[5]), .A2(cur_inst_addr_i[4]), .A3(
        cur_inst_addr_i[3]), .A4(cur_inst_addr_i[31]), .ZN(n244) );
  NOR4V0P5_8TH40 U356 ( .A1(cur_inst_addr_i[30]), .A2(cur_inst_addr_i[2]), 
        .A3(cur_inst_addr_i[29]), .A4(cur_inst_addr_i[28]), .ZN(n243) );
  NOR4V0P5_8TH40 U357 ( .A1(cur_inst_addr_i[27]), .A2(cur_inst_addr_i[26]), 
        .A3(cur_inst_addr_i[25]), .A4(cur_inst_addr_i[24]), .ZN(n242) );
  CLKNV1_8TH40 U358 ( .I(n248), .ZN(n247) );
  NOR2V0P5_8TH40 U359 ( .A1(n203), .A2(n28), .ZN(n246) );
  AOI221V0_8TH40 U360 ( .A1(n195), .A2(n252), .B1(n253), .B2(n28), .C(n248), 
        .ZN(n249) );
  OAI21V0_8TH40 U361 ( .A1(n136), .A2(n17), .B(n254), .ZN(n248) );
  AOAI211V0_8TH40 U362 ( .A1(n255), .A2(n39), .B(rst), .C(n251), .ZN(
        dmem_byte_sel[1]) );
  OAI31V0_8TH40 U363 ( .A1(n114), .A2(rst), .A3(n258), .B(n202), .ZN(n257) );
  NOR2V0P5_8TH40 U364 ( .A1(n195), .A2(n28), .ZN(n114) );
  CLKNV1_8TH40 U365 ( .I(n202), .ZN(n260) );
  CLKNAND2V1_8TH40 U366 ( .A1(n352), .A2(n261), .ZN(n202) );
  OAI211V0_8TH40 U367 ( .A1(n262), .A2(n39), .B(n255), .C(n258), .ZN(n259) );
  OA21V0_8TH40 U368 ( .A1(n28), .A2(n17), .B(n254), .Z(n255) );
  NOR2V0P5_8TH40 U369 ( .A1(n205), .A2(n264), .ZN(n263) );
  MUX2NV0_8TH40 U370 ( .I0(inst_type[3]), .I1(inst_type[0]), .S(inst_type[1]), 
        .ZN(n267) );
  CLKNV1_8TH40 U371 ( .I(n36), .ZN(n28) );
  NAND3V0P5_8TH40 U372 ( .A1(n268), .A2(n269), .A3(n209), .ZN(n252) );
  AND2V0_8TH40 U373 ( .A1(dmem_addr_i[9]), .A2(dmem_ce), .Z(dmem_addr_o[9]) );
  AND2V0_8TH40 U374 ( .A1(dmem_addr_i[8]), .A2(dmem_ce), .Z(dmem_addr_o[8]) );
  AND2V0_8TH40 U375 ( .A1(dmem_addr_i[7]), .A2(dmem_ce), .Z(dmem_addr_o[7]) );
  AND2V0_8TH40 U376 ( .A1(dmem_addr_i[6]), .A2(dmem_ce), .Z(dmem_addr_o[6]) );
  AND2V0_8TH40 U377 ( .A1(dmem_addr_i[5]), .A2(dmem_ce), .Z(dmem_addr_o[5]) );
  AND2V0_8TH40 U378 ( .A1(dmem_addr_i[4]), .A2(dmem_ce), .Z(dmem_addr_o[4]) );
  AND2V0_8TH40 U379 ( .A1(dmem_addr_i[3]), .A2(dmem_ce), .Z(dmem_addr_o[3]) );
  AND2V0_8TH40 U380 ( .A1(dmem_addr_i[31]), .A2(dmem_ce), .Z(dmem_addr_o[31])
         );
  AND2V0_8TH40 U381 ( .A1(dmem_addr_i[30]), .A2(dmem_ce), .Z(dmem_addr_o[30])
         );
  AND2V0_8TH40 U382 ( .A1(dmem_addr_i[2]), .A2(dmem_ce), .Z(dmem_addr_o[2]) );
  AND2V0_8TH40 U383 ( .A1(dmem_addr_i[29]), .A2(dmem_ce), .Z(dmem_addr_o[29])
         );
  AND2V0_8TH40 U384 ( .A1(dmem_addr_i[28]), .A2(dmem_ce), .Z(dmem_addr_o[28])
         );
  AND2V0_8TH40 U385 ( .A1(dmem_addr_i[27]), .A2(dmem_ce), .Z(dmem_addr_o[27])
         );
  AND2V0_8TH40 U386 ( .A1(dmem_addr_i[26]), .A2(dmem_ce), .Z(dmem_addr_o[26])
         );
  AND2V0_8TH40 U387 ( .A1(dmem_addr_i[25]), .A2(dmem_ce), .Z(dmem_addr_o[25])
         );
  AND2V0_8TH40 U388 ( .A1(dmem_addr_i[24]), .A2(dmem_ce), .Z(dmem_addr_o[24])
         );
  AND2V0_8TH40 U389 ( .A1(dmem_addr_i[23]), .A2(dmem_ce), .Z(dmem_addr_o[23])
         );
  AND2V0_8TH40 U390 ( .A1(dmem_addr_i[22]), .A2(dmem_ce), .Z(dmem_addr_o[22])
         );
  AND2V0_8TH40 U391 ( .A1(dmem_addr_i[21]), .A2(dmem_ce), .Z(dmem_addr_o[21])
         );
  AND2V0_8TH40 U392 ( .A1(dmem_addr_i[20]), .A2(dmem_ce), .Z(dmem_addr_o[20])
         );
  NOR2V0P5_8TH40 U393 ( .A1(n270), .A2(n271), .ZN(dmem_addr_o[1]) );
  AND2V0_8TH40 U394 ( .A1(dmem_addr_i[19]), .A2(dmem_ce), .Z(dmem_addr_o[19])
         );
  AND2V0_8TH40 U395 ( .A1(dmem_addr_i[18]), .A2(dmem_ce), .Z(dmem_addr_o[18])
         );
  AND2V0_8TH40 U396 ( .A1(dmem_addr_i[17]), .A2(dmem_ce), .Z(dmem_addr_o[17])
         );
  AND2V0_8TH40 U397 ( .A1(dmem_addr_i[16]), .A2(dmem_ce), .Z(dmem_addr_o[16])
         );
  AND2V0_8TH40 U398 ( .A1(dmem_addr_i[15]), .A2(dmem_ce), .Z(dmem_addr_o[15])
         );
  AND2V0_8TH40 U399 ( .A1(dmem_addr_i[14]), .A2(dmem_ce), .Z(dmem_addr_o[14])
         );
  AND2V0_8TH40 U400 ( .A1(dmem_addr_i[13]), .A2(dmem_ce), .Z(dmem_addr_o[13])
         );
  AND2V0_8TH40 U401 ( .A1(dmem_addr_i[12]), .A2(dmem_ce), .Z(dmem_addr_o[12])
         );
  AND2V0_8TH40 U402 ( .A1(dmem_addr_i[11]), .A2(dmem_ce), .Z(dmem_addr_o[11])
         );
  AND2V0_8TH40 U403 ( .A1(dmem_addr_i[10]), .A2(dmem_ce), .Z(dmem_addr_o[10])
         );
  OAI31V0_8TH40 U404 ( .A1(n194), .A2(n203), .A3(n204), .B(n1), .ZN(n272) );
  CLKNV1_8TH40 U405 ( .I(n115), .ZN(n194) );
  NAND3V0P5_8TH40 U406 ( .A1(n273), .A2(n274), .A3(inst_type[2]), .ZN(n115) );
  CLKNAND2V1_8TH40 U407 ( .A1(n153), .A2(n1), .ZN(n65) );
  CLKNV1_8TH40 U408 ( .I(n189), .ZN(n153) );
  NAND3V0P5_8TH40 U409 ( .A1(n266), .A2(n274), .A3(n273), .ZN(n189) );
  NOR2V0P5_8TH40 U410 ( .A1(n275), .A2(n271), .ZN(dmem_addr_o[0]) );
  CLKNV1_8TH40 U411 ( .I(n4), .ZN(n1) );
  CLKNAND2V1_8TH40 U412 ( .A1(n277), .A2(n352), .ZN(n4) );
  OAI31V0_8TH40 U413 ( .A1(n162), .A2(inst_type[3]), .A3(n278), .B(n3), .ZN(
        n40) );
  NAND3V0P5_8TH40 U414 ( .A1(n191), .A2(n274), .A3(inst_type[4]), .ZN(n3) );
  NAND3V0P5_8TH40 U415 ( .A1(n17), .A2(n207), .A3(n209), .ZN(n276) );
  INAND2V0_8TH40 U416 ( .A1(inst_type[0]), .B1(n279), .ZN(n209) );
  CLKNAND2V1_8TH40 U417 ( .A1(inst_type[0]), .A2(n279), .ZN(n17) );
  NOR3V0P5_8TH40 U418 ( .A1(inst_type[3]), .A2(inst_type[4]), .A3(inst_type[1]), .ZN(n279) );
  INOR2V0_8TH40 U419 ( .A1(cp0_we_i), .B1(rst), .ZN(cp0_we_o) );
  INOR2V0_8TH40 U420 ( .A1(cp0_wdata_i[9]), .B1(rst), .ZN(cp0_wdata_o[9]) );
  INOR2V0_8TH40 U421 ( .A1(cp0_wdata_i[8]), .B1(rst), .ZN(cp0_wdata_o[8]) );
  INOR2V0_8TH40 U422 ( .A1(cp0_wdata_i[7]), .B1(rst), .ZN(cp0_wdata_o[7]) );
  INOR2V0_8TH40 U423 ( .A1(cp0_wdata_i[6]), .B1(rst), .ZN(cp0_wdata_o[6]) );
  INOR2V0_8TH40 U424 ( .A1(cp0_wdata_i[5]), .B1(rst), .ZN(cp0_wdata_o[5]) );
  INOR2V0_8TH40 U425 ( .A1(cp0_wdata_i[4]), .B1(rst), .ZN(cp0_wdata_o[4]) );
  INOR2V0_8TH40 U426 ( .A1(cp0_wdata_i[3]), .B1(rst), .ZN(cp0_wdata_o[3]) );
  INOR2V0_8TH40 U427 ( .A1(cp0_wdata_i[31]), .B1(rst), .ZN(cp0_wdata_o[31]) );
  INOR2V0_8TH40 U428 ( .A1(cp0_wdata_i[30]), .B1(rst), .ZN(cp0_wdata_o[30]) );
  INOR2V0_8TH40 U429 ( .A1(cp0_wdata_i[2]), .B1(rst), .ZN(cp0_wdata_o[2]) );
  INOR2V0_8TH40 U430 ( .A1(cp0_wdata_i[29]), .B1(rst), .ZN(cp0_wdata_o[29]) );
  INOR2V0_8TH40 U431 ( .A1(cp0_wdata_i[28]), .B1(rst), .ZN(cp0_wdata_o[28]) );
  INOR2V0_8TH40 U432 ( .A1(cp0_wdata_i[27]), .B1(rst), .ZN(cp0_wdata_o[27]) );
  INOR2V0_8TH40 U433 ( .A1(cp0_wdata_i[26]), .B1(rst), .ZN(cp0_wdata_o[26]) );
  INOR2V0_8TH40 U434 ( .A1(cp0_wdata_i[25]), .B1(rst), .ZN(cp0_wdata_o[25]) );
  INOR2V0_8TH40 U435 ( .A1(cp0_wdata_i[24]), .B1(rst), .ZN(cp0_wdata_o[24]) );
  INOR2V0_8TH40 U436 ( .A1(cp0_wdata_i[23]), .B1(rst), .ZN(cp0_wdata_o[23]) );
  INOR2V0_8TH40 U437 ( .A1(cp0_wdata_i[22]), .B1(rst), .ZN(cp0_wdata_o[22]) );
  INOR2V0_8TH40 U438 ( .A1(cp0_wdata_i[21]), .B1(rst), .ZN(cp0_wdata_o[21]) );
  INOR2V0_8TH40 U439 ( .A1(cp0_wdata_i[20]), .B1(rst), .ZN(cp0_wdata_o[20]) );
  INOR2V0_8TH40 U440 ( .A1(cp0_wdata_i[1]), .B1(rst), .ZN(cp0_wdata_o[1]) );
  INOR2V0_8TH40 U441 ( .A1(cp0_wdata_i[19]), .B1(rst), .ZN(cp0_wdata_o[19]) );
  INOR2V0_8TH40 U442 ( .A1(cp0_wdata_i[18]), .B1(rst), .ZN(cp0_wdata_o[18]) );
  INOR2V0_8TH40 U443 ( .A1(cp0_wdata_i[17]), .B1(rst), .ZN(cp0_wdata_o[17]) );
  INOR2V0_8TH40 U444 ( .A1(cp0_wdata_i[16]), .B1(rst), .ZN(cp0_wdata_o[16]) );
  INOR2V0_8TH40 U445 ( .A1(cp0_wdata_i[15]), .B1(rst), .ZN(cp0_wdata_o[15]) );
  INOR2V0_8TH40 U446 ( .A1(cp0_wdata_i[14]), .B1(rst), .ZN(cp0_wdata_o[14]) );
  INOR2V0_8TH40 U447 ( .A1(cp0_wdata_i[13]), .B1(rst), .ZN(cp0_wdata_o[13]) );
  INOR2V0_8TH40 U448 ( .A1(cp0_wdata_i[12]), .B1(rst), .ZN(cp0_wdata_o[12]) );
  INOR2V0_8TH40 U449 ( .A1(cp0_wdata_i[11]), .B1(rst), .ZN(cp0_wdata_o[11]) );
  INOR2V0_8TH40 U450 ( .A1(cp0_wdata_i[10]), .B1(rst), .ZN(cp0_wdata_o[10]) );
  INOR2V0_8TH40 U451 ( .A1(cp0_wdata_i[0]), .B1(rst), .ZN(cp0_wdata_o[0]) );
  INOR2V0_8TH40 U452 ( .A1(cp0_waddr_i[4]), .B1(rst), .ZN(cp0_waddr_o[4]) );
  INOR2V0_8TH40 U453 ( .A1(cp0_waddr_i[3]), .B1(rst), .ZN(cp0_waddr_o[3]) );
  INOR2V0_8TH40 U454 ( .A1(cp0_waddr_i[2]), .B1(rst), .ZN(cp0_waddr_o[2]) );
  INOR2V0_8TH40 U455 ( .A1(cp0_waddr_i[1]), .B1(rst), .ZN(cp0_waddr_o[1]) );
  INOR2V0_8TH40 U456 ( .A1(cp0_waddr_i[0]), .B1(rst), .ZN(cp0_waddr_o[0]) );
  AO22V0_8TH40 U457 ( .A1(n280), .A2(wb_cp0_wdata[9]), .B1(cp0_epc_i[9]), .B2(
        n281), .Z(cp0_epc_o[9]) );
  AO22V0_8TH40 U458 ( .A1(n280), .A2(wb_cp0_wdata[8]), .B1(cp0_epc_i[8]), .B2(
        n281), .Z(cp0_epc_o[8]) );
  AO22V0_8TH40 U459 ( .A1(wb_cp0_wdata[7]), .A2(n280), .B1(cp0_epc_i[7]), .B2(
        n281), .Z(cp0_epc_o[7]) );
  AO22V0_8TH40 U460 ( .A1(wb_cp0_wdata[6]), .A2(n280), .B1(cp0_epc_i[6]), .B2(
        n281), .Z(cp0_epc_o[6]) );
  AO22V0_8TH40 U461 ( .A1(wb_cp0_wdata[5]), .A2(n280), .B1(cp0_epc_i[5]), .B2(
        n281), .Z(cp0_epc_o[5]) );
  AO22V0_8TH40 U462 ( .A1(wb_cp0_wdata[4]), .A2(n280), .B1(cp0_epc_i[4]), .B2(
        n281), .Z(cp0_epc_o[4]) );
  AO22V0_8TH40 U463 ( .A1(wb_cp0_wdata[3]), .A2(n280), .B1(cp0_epc_i[3]), .B2(
        n281), .Z(cp0_epc_o[3]) );
  AO22V0_8TH40 U464 ( .A1(wb_cp0_wdata[31]), .A2(n280), .B1(cp0_epc_i[31]), 
        .B2(n281), .Z(cp0_epc_o[31]) );
  AO22V0_8TH40 U465 ( .A1(wb_cp0_wdata[30]), .A2(n280), .B1(cp0_epc_i[30]), 
        .B2(n281), .Z(cp0_epc_o[30]) );
  AO22V0_8TH40 U466 ( .A1(wb_cp0_wdata[2]), .A2(n280), .B1(cp0_epc_i[2]), .B2(
        n281), .Z(cp0_epc_o[2]) );
  AO22V0_8TH40 U467 ( .A1(wb_cp0_wdata[29]), .A2(n280), .B1(cp0_epc_i[29]), 
        .B2(n281), .Z(cp0_epc_o[29]) );
  AO22V0_8TH40 U468 ( .A1(wb_cp0_wdata[28]), .A2(n280), .B1(cp0_epc_i[28]), 
        .B2(n281), .Z(cp0_epc_o[28]) );
  AO22V0_8TH40 U469 ( .A1(wb_cp0_wdata[27]), .A2(n280), .B1(cp0_epc_i[27]), 
        .B2(n281), .Z(cp0_epc_o[27]) );
  AO22V0_8TH40 U470 ( .A1(wb_cp0_wdata[26]), .A2(n280), .B1(cp0_epc_i[26]), 
        .B2(n281), .Z(cp0_epc_o[26]) );
  AO22V0_8TH40 U471 ( .A1(wb_cp0_wdata[25]), .A2(n280), .B1(cp0_epc_i[25]), 
        .B2(n281), .Z(cp0_epc_o[25]) );
  AO22V0_8TH40 U472 ( .A1(wb_cp0_wdata[24]), .A2(n280), .B1(cp0_epc_i[24]), 
        .B2(n281), .Z(cp0_epc_o[24]) );
  AO22V0_8TH40 U473 ( .A1(wb_cp0_wdata[23]), .A2(n280), .B1(cp0_epc_i[23]), 
        .B2(n281), .Z(cp0_epc_o[23]) );
  AO22V0_8TH40 U474 ( .A1(wb_cp0_wdata[22]), .A2(n280), .B1(cp0_epc_i[22]), 
        .B2(n281), .Z(cp0_epc_o[22]) );
  AO22V0_8TH40 U475 ( .A1(wb_cp0_wdata[21]), .A2(n280), .B1(cp0_epc_i[21]), 
        .B2(n281), .Z(cp0_epc_o[21]) );
  AO22V0_8TH40 U476 ( .A1(wb_cp0_wdata[20]), .A2(n280), .B1(cp0_epc_i[20]), 
        .B2(n281), .Z(cp0_epc_o[20]) );
  AO22V0_8TH40 U477 ( .A1(n280), .A2(wb_cp0_wdata[1]), .B1(cp0_epc_i[1]), .B2(
        n281), .Z(cp0_epc_o[1]) );
  AO22V0_8TH40 U478 ( .A1(wb_cp0_wdata[19]), .A2(n280), .B1(cp0_epc_i[19]), 
        .B2(n281), .Z(cp0_epc_o[19]) );
  AO22V0_8TH40 U479 ( .A1(wb_cp0_wdata[18]), .A2(n280), .B1(cp0_epc_i[18]), 
        .B2(n281), .Z(cp0_epc_o[18]) );
  AO22V0_8TH40 U480 ( .A1(wb_cp0_wdata[17]), .A2(n280), .B1(cp0_epc_i[17]), 
        .B2(n281), .Z(cp0_epc_o[17]) );
  AO22V0_8TH40 U481 ( .A1(wb_cp0_wdata[16]), .A2(n280), .B1(cp0_epc_i[16]), 
        .B2(n281), .Z(cp0_epc_o[16]) );
  AO22V0_8TH40 U482 ( .A1(n280), .A2(wb_cp0_wdata[15]), .B1(cp0_epc_i[15]), 
        .B2(n281), .Z(cp0_epc_o[15]) );
  AO22V0_8TH40 U483 ( .A1(n280), .A2(wb_cp0_wdata[14]), .B1(cp0_epc_i[14]), 
        .B2(n281), .Z(cp0_epc_o[14]) );
  AO22V0_8TH40 U484 ( .A1(n280), .A2(wb_cp0_wdata[13]), .B1(cp0_epc_i[13]), 
        .B2(n281), .Z(cp0_epc_o[13]) );
  AO22V0_8TH40 U485 ( .A1(n280), .A2(wb_cp0_wdata[12]), .B1(cp0_epc_i[12]), 
        .B2(n281), .Z(cp0_epc_o[12]) );
  AO22V0_8TH40 U486 ( .A1(n280), .A2(wb_cp0_wdata[11]), .B1(cp0_epc_i[11]), 
        .B2(n281), .Z(cp0_epc_o[11]) );
  AO22V0_8TH40 U487 ( .A1(n280), .A2(wb_cp0_wdata[10]), .B1(cp0_epc_i[10]), 
        .B2(n281), .Z(cp0_epc_o[10]) );
  AO22V0_8TH40 U488 ( .A1(wb_cp0_wdata[0]), .A2(n280), .B1(cp0_epc_i[0]), .B2(
        n281), .Z(cp0_epc_o[0]) );
  INOR2V0_8TH40 U489 ( .A1(n282), .B1(rst), .ZN(n281) );
  NOR2V0P5_8TH40 U490 ( .A1(n282), .A2(rst), .ZN(n280) );
  I2NAND3V1_8TH40 U491 ( .A1(wb_cp0_waddr[0]), .A2(n233), .B(wb_cp0_waddr[1]), 
        .ZN(n282) );
  INAND4V0_8TH40 U492 ( .A1(wb_cp0_waddr[4]), .B1(wb_cp0_waddr[2]), .B2(
        wb_cp0_we), .B3(wb_cp0_waddr[3]), .ZN(n233) );
  AOI22V0_8TH40 U493 ( .A1(n287), .A2(ls_data_tmp[7]), .B1(n288), .B2(
        ls_data_tmp[15]), .ZN(n286) );
  AOI22V0_8TH40 U494 ( .A1(n287), .A2(ls_data_tmp[6]), .B1(n288), .B2(
        ls_data_tmp[14]), .ZN(n290) );
  AOI22V0_8TH40 U495 ( .A1(n287), .A2(ls_data_tmp[5]), .B1(n288), .B2(
        ls_data_tmp[13]), .ZN(n292) );
  AOI22V0_8TH40 U496 ( .A1(n287), .A2(ls_data_tmp[4]), .B1(n288), .B2(
        ls_data_tmp[12]), .ZN(n294) );
  AOI22V0_8TH40 U497 ( .A1(n287), .A2(ls_data_tmp[3]), .B1(n288), .B2(
        ls_data_tmp[11]), .ZN(n296) );
  AOI22V0_8TH40 U498 ( .A1(n287), .A2(ls_data_tmp[2]), .B1(n288), .B2(
        ls_data_tmp[10]), .ZN(n298) );
  AOI22V0_8TH40 U499 ( .A1(n287), .A2(ls_data_tmp[1]), .B1(n288), .B2(
        ls_data_tmp[9]), .ZN(n300) );
  AOI22V0_8TH40 U500 ( .A1(n287), .A2(ls_data_tmp[0]), .B1(n288), .B2(
        ls_data_tmp[8]), .ZN(n302) );
  OAOI211V0_8TH40 U501 ( .A1(n269), .A2(n188), .B(n262), .C(rst), .ZN(n288) );
  OAOI211V0_8TH40 U502 ( .A1(n269), .A2(n36), .B(n268), .C(rst), .ZN(n287) );
  AOI22V0_8TH40 U503 ( .A1(n305), .A2(ls_data_tmp[7]), .B1(n306), .B2(
        ls_data_tmp[23]), .ZN(n304) );
  CLKNV1_8TH40 U504 ( .I(ls_data_tmp[31]), .ZN(n283) );
  AOI22V0_8TH40 U505 ( .A1(n305), .A2(ls_data_tmp[6]), .B1(n306), .B2(
        ls_data_tmp[22]), .ZN(n307) );
  CLKNV1_8TH40 U506 ( .I(ls_data_tmp[30]), .ZN(n73) );
  AOI22V0_8TH40 U507 ( .A1(n305), .A2(ls_data_tmp[5]), .B1(n306), .B2(
        ls_data_tmp[21]), .ZN(n308) );
  CLKNV1_8TH40 U508 ( .I(ls_data_tmp[29]), .ZN(n84) );
  AOI22V0_8TH40 U509 ( .A1(n305), .A2(ls_data_tmp[4]), .B1(n306), .B2(
        ls_data_tmp[20]), .ZN(n309) );
  CLKNV1_8TH40 U510 ( .I(ls_data_tmp[28]), .ZN(n90) );
  AOI22V0_8TH40 U511 ( .A1(n305), .A2(ls_data_tmp[3]), .B1(n306), .B2(
        ls_data_tmp[19]), .ZN(n310) );
  CLKNV1_8TH40 U512 ( .I(ls_data_tmp[27]), .ZN(n96) );
  AOI22V0_8TH40 U513 ( .A1(n305), .A2(ls_data_tmp[2]), .B1(n306), .B2(
        ls_data_tmp[18]), .ZN(n311) );
  CLKNV1_8TH40 U514 ( .I(ls_data_tmp[26]), .ZN(n102) );
  AOI22V0_8TH40 U515 ( .A1(n305), .A2(ls_data_tmp[1]), .B1(n306), .B2(
        ls_data_tmp[17]), .ZN(n312) );
  CLKNV1_8TH40 U516 ( .I(ls_data_tmp[25]), .ZN(n108) );
  AOI22V0_8TH40 U517 ( .A1(n305), .A2(ls_data_tmp[0]), .B1(n306), .B2(
        ls_data_tmp[16]), .ZN(n313) );
  CLKNV1_8TH40 U518 ( .I(n284), .ZN(n306) );
  OAI21V0_8TH40 U519 ( .A1(n264), .A2(n314), .B(n352), .ZN(n284) );
  CLKNAND2V1_8TH40 U520 ( .A1(n195), .A2(n203), .ZN(n315) );
  CLKNV1_8TH40 U521 ( .I(ls_data_tmp[24]), .ZN(n113) );
  AOI22V0_8TH40 U522 ( .A1(n320), .A2(ls_data_tmp[23]), .B1(n321), .B2(
        ls_data_tmp[31]), .ZN(n319) );
  CLKNV1_8TH40 U523 ( .I(ls_data_tmp[7]), .ZN(n317) );
  AOI22V0_8TH40 U524 ( .A1(n320), .A2(ls_data_tmp[22]), .B1(n321), .B2(
        ls_data_tmp[30]), .ZN(n323) );
  CLKNV1_8TH40 U525 ( .I(ls_data_tmp[6]), .ZN(n322) );
  AOI22V0_8TH40 U526 ( .A1(n320), .A2(ls_data_tmp[21]), .B1(n321), .B2(
        ls_data_tmp[29]), .ZN(n325) );
  CLKNV1_8TH40 U527 ( .I(ls_data_tmp[5]), .ZN(n324) );
  AOI22V0_8TH40 U528 ( .A1(n320), .A2(ls_data_tmp[20]), .B1(n321), .B2(
        ls_data_tmp[28]), .ZN(n327) );
  CLKNV1_8TH40 U529 ( .I(ls_data_tmp[4]), .ZN(n326) );
  AOI22V0_8TH40 U530 ( .A1(n320), .A2(ls_data_tmp[19]), .B1(n321), .B2(
        ls_data_tmp[27]), .ZN(n329) );
  CLKNV1_8TH40 U531 ( .I(ls_data_tmp[3]), .ZN(n328) );
  AOI22V0_8TH40 U532 ( .A1(n320), .A2(ls_data_tmp[18]), .B1(n321), .B2(
        ls_data_tmp[26]), .ZN(n331) );
  CLKNV1_8TH40 U533 ( .I(ls_data_tmp[2]), .ZN(n330) );
  AOI22V0_8TH40 U534 ( .A1(n320), .A2(ls_data_tmp[17]), .B1(n321), .B2(
        ls_data_tmp[25]), .ZN(n334) );
  CLKNV1_8TH40 U535 ( .I(ls_data_tmp[1]), .ZN(n332) );
  AOI22V0_8TH40 U536 ( .A1(n320), .A2(ls_data_tmp[16]), .B1(n321), .B2(
        ls_data_tmp[24]), .ZN(n336) );
  CLKNV1_8TH40 U537 ( .I(n337), .ZN(n321) );
  CLKNV1_8TH40 U538 ( .I(n303), .ZN(n320) );
  CLKNV1_8TH40 U539 ( .I(ls_data_tmp[0]), .ZN(n335) );
  OA21V0_8TH40 U540 ( .A1(rst), .A2(n268), .B(n250), .Z(n316) );
  NAND3V0P5_8TH40 U541 ( .A1(n136), .A2(n352), .A3(n203), .ZN(n250) );
  CLKNV1_8TH40 U542 ( .I(n269), .ZN(n203) );
  AOI22V0_8TH40 U543 ( .A1(ls_data_tmp[7]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[31]), .ZN(n338) );
  CLKNV1_8TH40 U544 ( .I(ls_data_tmp[23]), .ZN(n285) );
  CLKNV1_8TH40 U545 ( .I(ls_data_tmp[15]), .ZN(n163) );
  AOI22V0_8TH40 U546 ( .A1(ls_data_tmp[6]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[30]), .ZN(n341) );
  CLKNV1_8TH40 U547 ( .I(ls_data_tmp[22]), .ZN(n289) );
  CLKNV1_8TH40 U548 ( .I(ls_data_tmp[14]), .ZN(n169) );
  AOI22V0_8TH40 U549 ( .A1(ls_data_tmp[5]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[29]), .ZN(n342) );
  CLKNV1_8TH40 U550 ( .I(ls_data_tmp[21]), .ZN(n291) );
  CLKNV1_8TH40 U551 ( .I(ls_data_tmp[13]), .ZN(n174) );
  AOI22V0_8TH40 U552 ( .A1(ls_data_tmp[4]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[28]), .ZN(n343) );
  CLKNV1_8TH40 U553 ( .I(ls_data_tmp[20]), .ZN(n293) );
  CLKNV1_8TH40 U554 ( .I(ls_data_tmp[12]), .ZN(n179) );
  AOI22V0_8TH40 U555 ( .A1(ls_data_tmp[3]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[27]), .ZN(n344) );
  CLKNV1_8TH40 U556 ( .I(ls_data_tmp[19]), .ZN(n295) );
  CLKNV1_8TH40 U557 ( .I(ls_data_tmp[11]), .ZN(n184) );
  AOI22V0_8TH40 U558 ( .A1(ls_data_tmp[2]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[26]), .ZN(n345) );
  CLKNV1_8TH40 U559 ( .I(ls_data_tmp[18]), .ZN(n297) );
  CLKNV1_8TH40 U560 ( .I(ls_data_tmp[10]), .ZN(n193) );
  AOI22V0_8TH40 U561 ( .A1(ls_data_tmp[1]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[25]), .ZN(n346) );
  CLKNV1_8TH40 U562 ( .I(ls_data_tmp[17]), .ZN(n299) );
  CLKNV1_8TH40 U563 ( .I(ls_data_tmp[9]), .ZN(n15) );
  AOI22V0_8TH40 U564 ( .A1(ls_data_tmp[0]), .A2(n339), .B1(n340), .B2(
        ls_data_tmp[24]), .ZN(n347) );
  INOR2V0_8TH40 U565 ( .A1(n256), .B1(n258), .ZN(n340) );
  NOR2V0P5_8TH40 U566 ( .A1(n192), .A2(rst), .ZN(n256) );
  OAI21V0_8TH40 U567 ( .A1(rst), .A2(n268), .B(n318), .ZN(n339) );
  OAI31V0_8TH40 U568 ( .A1(n314), .A2(n253), .A3(n264), .B(n352), .ZN(n318) );
  CLKNAND2V1_8TH40 U569 ( .A1(n348), .A2(n349), .ZN(n264) );
  OAI22V0_8TH40 U570 ( .A1(n192), .A2(n269), .B1(n36), .B2(n258), .ZN(n314) );
  CLKNAND2V1_8TH40 U571 ( .A1(n270), .A2(n275), .ZN(n36) );
  CLKNAND2V1_8TH40 U572 ( .A1(dmem_addr_i[0]), .A2(dmem_addr_i[1]), .ZN(n192)
         );
  NAND3V0P5_8TH40 U573 ( .A1(n136), .A2(n352), .A3(n204), .ZN(n337) );
  CLKNV1_8TH40 U574 ( .I(n39), .ZN(n136) );
  CLKNAND2V1_8TH40 U575 ( .A1(dmem_addr_i[1]), .A2(n275), .ZN(n39) );
  CLKNV1_8TH40 U576 ( .I(dmem_addr_i[0]), .ZN(n275) );
  CLKNV1_8TH40 U577 ( .I(ls_data_tmp[16]), .ZN(n301) );
  NAND3V0P5_8TH40 U578 ( .A1(n195), .A2(n352), .A3(n204), .ZN(n303) );
  CLKNV1_8TH40 U579 ( .I(n188), .ZN(n195) );
  CLKNAND2V1_8TH40 U580 ( .A1(dmem_addr_i[0]), .A2(n270), .ZN(n188) );
  CLKNV1_8TH40 U581 ( .I(dmem_addr_i[1]), .ZN(n270) );
  CLKNV1_8TH40 U582 ( .I(ls_data_tmp[8]), .ZN(n25) );
  CLKNAND2V1_8TH40 U583 ( .A1(n352), .A2(n217), .ZN(N569) );
  CLKNV1_8TH40 U584 ( .I(n261), .ZN(n277) );
  NAND3V0P5_8TH40 U585 ( .A1(inst_type[6]), .A2(inst_type[5]), .A3(
        inst_type[7]), .ZN(n261) );
  NAND3V0P5_8TH40 U586 ( .A1(n262), .A2(n268), .A3(n349), .ZN(n206) );
  I2NAND3V1_8TH40 U587 ( .A1(n162), .A2(n278), .B(inst_type[3]), .ZN(n349) );
  NAND3V0P5_8TH40 U588 ( .A1(n191), .A2(n265), .A3(inst_type[3]), .ZN(n268) );
  CLKNV1_8TH40 U589 ( .I(n253), .ZN(n262) );
  NOR3V0P5_8TH40 U590 ( .A1(n274), .A2(inst_type[1]), .A3(n162), .ZN(n253) );
  NAND3V0P5_8TH40 U591 ( .A1(n266), .A2(n265), .A3(inst_type[0]), .ZN(n162) );
  CLKNV1_8TH40 U592 ( .I(inst_type[4]), .ZN(n265) );
  CLKNV1_8TH40 U593 ( .I(inst_type[3]), .ZN(n274) );
  CLKNV1_8TH40 U594 ( .I(n258), .ZN(n204) );
  NAND3V0P5_8TH40 U595 ( .A1(inst_type[3]), .A2(n266), .A3(n273), .ZN(n258) );
  CLKNV1_8TH40 U596 ( .I(inst_type[2]), .ZN(n266) );
  CLKNAND2V1_8TH40 U597 ( .A1(n269), .A2(n207), .ZN(n350) );
  CKMUX2V2_8TH40 U598 ( .I0(llbit_i), .I1(wb_llbit_value), .S(wb_llbit_we), 
        .Z(n351) );
  NAND3V0P5_8TH40 U599 ( .A1(inst_type[3]), .A2(n191), .A3(inst_type[4]), .ZN(
        n348) );
  NOR3V0P5_8TH40 U600 ( .A1(inst_type[1]), .A2(inst_type[2]), .A3(inst_type[0]), .ZN(n191) );
  NAND3V0P5_8TH40 U601 ( .A1(n273), .A2(inst_type[3]), .A3(inst_type[2]), .ZN(
        n269) );
  NOR3V0P5_8TH40 U602 ( .A1(inst_type[0]), .A2(inst_type[4]), .A3(n278), .ZN(
        n273) );
  CLKNV1_8TH40 U603 ( .I(inst_type[1]), .ZN(n278) );
  CLKNV1_8TH40 U604 ( .I(rst), .ZN(n352) );
endmodule


module pipe_reg_memwb ( clk, rst, stall_ctrl, mem_gpr_we, mem_target_gpr, 
        mem_exe_result, mem_hi, mem_lo, mem_hilo_we, mem_llbit_we, 
        mem_llbit_value, mem_cp0_we, mem_cp0_waddr, mem_cp0_wdata, wb_gpr_we, 
        wb_target_gpr, wb_exe_result, wb_hi, wb_lo, wb_hilo_we, wb_llbit_we, 
        wb_llbit_value, wb_cp0_we, wb_cp0_waddr, wb_cp0_wdata, flush_BAR );
  input [5:0] stall_ctrl;
  input [4:0] mem_target_gpr;
  input [31:0] mem_exe_result;
  input [31:0] mem_hi;
  input [31:0] mem_lo;
  input [4:0] mem_cp0_waddr;
  input [31:0] mem_cp0_wdata;
  output [4:0] wb_target_gpr;
  output [31:0] wb_exe_result;
  output [31:0] wb_hi;
  output [31:0] wb_lo;
  output [4:0] wb_cp0_waddr;
  output [31:0] wb_cp0_wdata;
  input clk, rst, mem_gpr_we, mem_hilo_we, mem_llbit_we, mem_llbit_value,
         mem_cp0_we, flush_BAR;
  output wb_gpr_we, wb_hilo_we, wb_llbit_we, wb_llbit_value, wb_cp0_we;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144;

  DQV4_8TH40 wb_cp0_we_reg ( .D(n144), .CK(clk), .Q(wb_cp0_we) );
  DQV4_8TH40 wb_cp0_waddr_reg_4_ ( .D(n143), .CK(clk), .Q(wb_cp0_waddr[4]) );
  DQV4_8TH40 wb_cp0_waddr_reg_3_ ( .D(n142), .CK(clk), .Q(wb_cp0_waddr[3]) );
  DQV4_8TH40 wb_cp0_waddr_reg_2_ ( .D(n141), .CK(clk), .Q(wb_cp0_waddr[2]) );
  DQV4_8TH40 wb_cp0_waddr_reg_1_ ( .D(n140), .CK(clk), .Q(wb_cp0_waddr[1]) );
  DQV4_8TH40 wb_cp0_waddr_reg_0_ ( .D(n139), .CK(clk), .Q(wb_cp0_waddr[0]) );
  DQV4_8TH40 wb_cp0_wdata_reg_31_ ( .D(n138), .CK(clk), .Q(wb_cp0_wdata[31])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_30_ ( .D(n137), .CK(clk), .Q(wb_cp0_wdata[30])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_29_ ( .D(n136), .CK(clk), .Q(wb_cp0_wdata[29])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_28_ ( .D(n135), .CK(clk), .Q(wb_cp0_wdata[28])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_27_ ( .D(n134), .CK(clk), .Q(wb_cp0_wdata[27])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_26_ ( .D(n133), .CK(clk), .Q(wb_cp0_wdata[26])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_25_ ( .D(n132), .CK(clk), .Q(wb_cp0_wdata[25])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_24_ ( .D(n131), .CK(clk), .Q(wb_cp0_wdata[24])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_23_ ( .D(n130), .CK(clk), .Q(wb_cp0_wdata[23])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_22_ ( .D(n129), .CK(clk), .Q(wb_cp0_wdata[22])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_21_ ( .D(n128), .CK(clk), .Q(wb_cp0_wdata[21])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_20_ ( .D(n127), .CK(clk), .Q(wb_cp0_wdata[20])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_19_ ( .D(n126), .CK(clk), .Q(wb_cp0_wdata[19])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_18_ ( .D(n125), .CK(clk), .Q(wb_cp0_wdata[18])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_17_ ( .D(n124), .CK(clk), .Q(wb_cp0_wdata[17])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_16_ ( .D(n123), .CK(clk), .Q(wb_cp0_wdata[16])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_15_ ( .D(n122), .CK(clk), .Q(wb_cp0_wdata[15])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_14_ ( .D(n121), .CK(clk), .Q(wb_cp0_wdata[14])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_13_ ( .D(n120), .CK(clk), .Q(wb_cp0_wdata[13])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_12_ ( .D(n119), .CK(clk), .Q(wb_cp0_wdata[12])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_11_ ( .D(n118), .CK(clk), .Q(wb_cp0_wdata[11])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_10_ ( .D(n117), .CK(clk), .Q(wb_cp0_wdata[10])
         );
  DQV4_8TH40 wb_cp0_wdata_reg_9_ ( .D(n116), .CK(clk), .Q(wb_cp0_wdata[9]) );
  DQV4_8TH40 wb_cp0_wdata_reg_8_ ( .D(n115), .CK(clk), .Q(wb_cp0_wdata[8]) );
  DQV4_8TH40 wb_cp0_wdata_reg_7_ ( .D(n114), .CK(clk), .Q(wb_cp0_wdata[7]) );
  DQV4_8TH40 wb_cp0_wdata_reg_6_ ( .D(n113), .CK(clk), .Q(wb_cp0_wdata[6]) );
  DQV4_8TH40 wb_cp0_wdata_reg_5_ ( .D(n112), .CK(clk), .Q(wb_cp0_wdata[5]) );
  DQV4_8TH40 wb_cp0_wdata_reg_4_ ( .D(n111), .CK(clk), .Q(wb_cp0_wdata[4]) );
  DQV4_8TH40 wb_cp0_wdata_reg_3_ ( .D(n110), .CK(clk), .Q(wb_cp0_wdata[3]) );
  DQV4_8TH40 wb_cp0_wdata_reg_2_ ( .D(n109), .CK(clk), .Q(wb_cp0_wdata[2]) );
  DQV4_8TH40 wb_cp0_wdata_reg_1_ ( .D(n108), .CK(clk), .Q(wb_cp0_wdata[1]) );
  DQV4_8TH40 wb_cp0_wdata_reg_0_ ( .D(n107), .CK(clk), .Q(wb_cp0_wdata[0]) );
  DQV4_8TH40 wb_gpr_we_reg ( .D(n106), .CK(clk), .Q(wb_gpr_we) );
  DQV4_8TH40 wb_target_gpr_reg_4_ ( .D(n105), .CK(clk), .Q(wb_target_gpr[4])
         );
  DQV4_8TH40 wb_target_gpr_reg_3_ ( .D(n104), .CK(clk), .Q(wb_target_gpr[3])
         );
  DQV4_8TH40 wb_target_gpr_reg_2_ ( .D(n103), .CK(clk), .Q(wb_target_gpr[2])
         );
  DQV4_8TH40 wb_target_gpr_reg_1_ ( .D(n102), .CK(clk), .Q(wb_target_gpr[1])
         );
  DQV4_8TH40 wb_target_gpr_reg_0_ ( .D(n101), .CK(clk), .Q(wb_target_gpr[0])
         );
  DQV4_8TH40 wb_exe_result_reg_31_ ( .D(n100), .CK(clk), .Q(wb_exe_result[31])
         );
  DQV4_8TH40 wb_exe_result_reg_30_ ( .D(n99), .CK(clk), .Q(wb_exe_result[30])
         );
  DQV4_8TH40 wb_exe_result_reg_29_ ( .D(n98), .CK(clk), .Q(wb_exe_result[29])
         );
  DQV4_8TH40 wb_exe_result_reg_28_ ( .D(n97), .CK(clk), .Q(wb_exe_result[28])
         );
  DQV4_8TH40 wb_exe_result_reg_27_ ( .D(n96), .CK(clk), .Q(wb_exe_result[27])
         );
  DQV4_8TH40 wb_exe_result_reg_26_ ( .D(n95), .CK(clk), .Q(wb_exe_result[26])
         );
  DQV4_8TH40 wb_exe_result_reg_25_ ( .D(n94), .CK(clk), .Q(wb_exe_result[25])
         );
  DQV4_8TH40 wb_exe_result_reg_24_ ( .D(n93), .CK(clk), .Q(wb_exe_result[24])
         );
  DQV4_8TH40 wb_exe_result_reg_23_ ( .D(n92), .CK(clk), .Q(wb_exe_result[23])
         );
  DQV4_8TH40 wb_exe_result_reg_22_ ( .D(n91), .CK(clk), .Q(wb_exe_result[22])
         );
  DQV4_8TH40 wb_exe_result_reg_21_ ( .D(n90), .CK(clk), .Q(wb_exe_result[21])
         );
  DQV4_8TH40 wb_exe_result_reg_20_ ( .D(n89), .CK(clk), .Q(wb_exe_result[20])
         );
  DQV4_8TH40 wb_exe_result_reg_19_ ( .D(n88), .CK(clk), .Q(wb_exe_result[19])
         );
  DQV4_8TH40 wb_exe_result_reg_18_ ( .D(n87), .CK(clk), .Q(wb_exe_result[18])
         );
  DQV4_8TH40 wb_exe_result_reg_17_ ( .D(n86), .CK(clk), .Q(wb_exe_result[17])
         );
  DQV4_8TH40 wb_exe_result_reg_16_ ( .D(n85), .CK(clk), .Q(wb_exe_result[16])
         );
  DQV4_8TH40 wb_exe_result_reg_15_ ( .D(n84), .CK(clk), .Q(wb_exe_result[15])
         );
  DQV4_8TH40 wb_exe_result_reg_14_ ( .D(n83), .CK(clk), .Q(wb_exe_result[14])
         );
  DQV4_8TH40 wb_exe_result_reg_13_ ( .D(n82), .CK(clk), .Q(wb_exe_result[13])
         );
  DQV4_8TH40 wb_exe_result_reg_12_ ( .D(n81), .CK(clk), .Q(wb_exe_result[12])
         );
  DQV4_8TH40 wb_exe_result_reg_11_ ( .D(n80), .CK(clk), .Q(wb_exe_result[11])
         );
  DQV4_8TH40 wb_exe_result_reg_10_ ( .D(n79), .CK(clk), .Q(wb_exe_result[10])
         );
  DQV4_8TH40 wb_exe_result_reg_9_ ( .D(n78), .CK(clk), .Q(wb_exe_result[9]) );
  DQV4_8TH40 wb_exe_result_reg_8_ ( .D(n77), .CK(clk), .Q(wb_exe_result[8]) );
  DQV4_8TH40 wb_exe_result_reg_7_ ( .D(n76), .CK(clk), .Q(wb_exe_result[7]) );
  DQV4_8TH40 wb_exe_result_reg_6_ ( .D(n75), .CK(clk), .Q(wb_exe_result[6]) );
  DQV4_8TH40 wb_exe_result_reg_5_ ( .D(n74), .CK(clk), .Q(wb_exe_result[5]) );
  DQV4_8TH40 wb_exe_result_reg_4_ ( .D(n73), .CK(clk), .Q(wb_exe_result[4]) );
  DQV4_8TH40 wb_exe_result_reg_3_ ( .D(n72), .CK(clk), .Q(wb_exe_result[3]) );
  DQV4_8TH40 wb_exe_result_reg_2_ ( .D(n71), .CK(clk), .Q(wb_exe_result[2]) );
  DQV4_8TH40 wb_exe_result_reg_1_ ( .D(n70), .CK(clk), .Q(wb_exe_result[1]) );
  DQV4_8TH40 wb_exe_result_reg_0_ ( .D(n69), .CK(clk), .Q(wb_exe_result[0]) );
  DQV4_8TH40 wb_hi_reg_31_ ( .D(n68), .CK(clk), .Q(wb_hi[31]) );
  DQV4_8TH40 wb_hi_reg_30_ ( .D(n67), .CK(clk), .Q(wb_hi[30]) );
  DQV4_8TH40 wb_hi_reg_29_ ( .D(n66), .CK(clk), .Q(wb_hi[29]) );
  DQV4_8TH40 wb_hi_reg_28_ ( .D(n65), .CK(clk), .Q(wb_hi[28]) );
  DQV4_8TH40 wb_hi_reg_27_ ( .D(n64), .CK(clk), .Q(wb_hi[27]) );
  DQV4_8TH40 wb_hi_reg_26_ ( .D(n63), .CK(clk), .Q(wb_hi[26]) );
  DQV4_8TH40 wb_hi_reg_25_ ( .D(n62), .CK(clk), .Q(wb_hi[25]) );
  DQV4_8TH40 wb_hi_reg_24_ ( .D(n61), .CK(clk), .Q(wb_hi[24]) );
  DQV4_8TH40 wb_hi_reg_23_ ( .D(n60), .CK(clk), .Q(wb_hi[23]) );
  DQV4_8TH40 wb_hi_reg_22_ ( .D(n59), .CK(clk), .Q(wb_hi[22]) );
  DQV4_8TH40 wb_hi_reg_21_ ( .D(n58), .CK(clk), .Q(wb_hi[21]) );
  DQV4_8TH40 wb_hi_reg_20_ ( .D(n57), .CK(clk), .Q(wb_hi[20]) );
  DQV4_8TH40 wb_hi_reg_19_ ( .D(n56), .CK(clk), .Q(wb_hi[19]) );
  DQV4_8TH40 wb_hi_reg_18_ ( .D(n55), .CK(clk), .Q(wb_hi[18]) );
  DQV4_8TH40 wb_hi_reg_17_ ( .D(n54), .CK(clk), .Q(wb_hi[17]) );
  DQV4_8TH40 wb_hi_reg_16_ ( .D(n53), .CK(clk), .Q(wb_hi[16]) );
  DQV4_8TH40 wb_hi_reg_15_ ( .D(n52), .CK(clk), .Q(wb_hi[15]) );
  DQV4_8TH40 wb_hi_reg_14_ ( .D(n51), .CK(clk), .Q(wb_hi[14]) );
  DQV4_8TH40 wb_hi_reg_13_ ( .D(n50), .CK(clk), .Q(wb_hi[13]) );
  DQV4_8TH40 wb_hi_reg_12_ ( .D(n49), .CK(clk), .Q(wb_hi[12]) );
  DQV4_8TH40 wb_hi_reg_11_ ( .D(n48), .CK(clk), .Q(wb_hi[11]) );
  DQV4_8TH40 wb_hi_reg_10_ ( .D(n47), .CK(clk), .Q(wb_hi[10]) );
  DQV4_8TH40 wb_hi_reg_9_ ( .D(n46), .CK(clk), .Q(wb_hi[9]) );
  DQV4_8TH40 wb_hi_reg_8_ ( .D(n45), .CK(clk), .Q(wb_hi[8]) );
  DQV4_8TH40 wb_hi_reg_7_ ( .D(n44), .CK(clk), .Q(wb_hi[7]) );
  DQV4_8TH40 wb_hi_reg_6_ ( .D(n43), .CK(clk), .Q(wb_hi[6]) );
  DQV4_8TH40 wb_hi_reg_5_ ( .D(n42), .CK(clk), .Q(wb_hi[5]) );
  DQV4_8TH40 wb_hi_reg_4_ ( .D(n41), .CK(clk), .Q(wb_hi[4]) );
  DQV4_8TH40 wb_hi_reg_3_ ( .D(n40), .CK(clk), .Q(wb_hi[3]) );
  DQV4_8TH40 wb_hi_reg_2_ ( .D(n39), .CK(clk), .Q(wb_hi[2]) );
  DQV4_8TH40 wb_hi_reg_1_ ( .D(n38), .CK(clk), .Q(wb_hi[1]) );
  DQV4_8TH40 wb_hi_reg_0_ ( .D(n37), .CK(clk), .Q(wb_hi[0]) );
  DQV4_8TH40 wb_lo_reg_31_ ( .D(n36), .CK(clk), .Q(wb_lo[31]) );
  DQV4_8TH40 wb_lo_reg_30_ ( .D(n35), .CK(clk), .Q(wb_lo[30]) );
  DQV4_8TH40 wb_lo_reg_29_ ( .D(n34), .CK(clk), .Q(wb_lo[29]) );
  DQV4_8TH40 wb_lo_reg_28_ ( .D(n33), .CK(clk), .Q(wb_lo[28]) );
  DQV4_8TH40 wb_lo_reg_27_ ( .D(n32), .CK(clk), .Q(wb_lo[27]) );
  DQV4_8TH40 wb_lo_reg_26_ ( .D(n31), .CK(clk), .Q(wb_lo[26]) );
  DQV4_8TH40 wb_lo_reg_25_ ( .D(n30), .CK(clk), .Q(wb_lo[25]) );
  DQV4_8TH40 wb_lo_reg_24_ ( .D(n29), .CK(clk), .Q(wb_lo[24]) );
  DQV4_8TH40 wb_lo_reg_23_ ( .D(n28), .CK(clk), .Q(wb_lo[23]) );
  DQV4_8TH40 wb_lo_reg_22_ ( .D(n27), .CK(clk), .Q(wb_lo[22]) );
  DQV4_8TH40 wb_lo_reg_21_ ( .D(n26), .CK(clk), .Q(wb_lo[21]) );
  DQV4_8TH40 wb_lo_reg_20_ ( .D(n25), .CK(clk), .Q(wb_lo[20]) );
  DQV4_8TH40 wb_lo_reg_19_ ( .D(n24), .CK(clk), .Q(wb_lo[19]) );
  DQV4_8TH40 wb_lo_reg_18_ ( .D(n23), .CK(clk), .Q(wb_lo[18]) );
  DQV4_8TH40 wb_lo_reg_17_ ( .D(n22), .CK(clk), .Q(wb_lo[17]) );
  DQV4_8TH40 wb_lo_reg_16_ ( .D(n21), .CK(clk), .Q(wb_lo[16]) );
  DQV4_8TH40 wb_lo_reg_15_ ( .D(n20), .CK(clk), .Q(wb_lo[15]) );
  DQV4_8TH40 wb_lo_reg_14_ ( .D(n19), .CK(clk), .Q(wb_lo[14]) );
  DQV4_8TH40 wb_lo_reg_13_ ( .D(n18), .CK(clk), .Q(wb_lo[13]) );
  DQV4_8TH40 wb_lo_reg_12_ ( .D(n17), .CK(clk), .Q(wb_lo[12]) );
  DQV4_8TH40 wb_lo_reg_11_ ( .D(n16), .CK(clk), .Q(wb_lo[11]) );
  DQV4_8TH40 wb_lo_reg_10_ ( .D(n15), .CK(clk), .Q(wb_lo[10]) );
  DQV4_8TH40 wb_lo_reg_9_ ( .D(n14), .CK(clk), .Q(wb_lo[9]) );
  DQV4_8TH40 wb_lo_reg_8_ ( .D(n13), .CK(clk), .Q(wb_lo[8]) );
  DQV4_8TH40 wb_lo_reg_7_ ( .D(n12), .CK(clk), .Q(wb_lo[7]) );
  DQV4_8TH40 wb_lo_reg_6_ ( .D(n11), .CK(clk), .Q(wb_lo[6]) );
  DQV4_8TH40 wb_lo_reg_5_ ( .D(n10), .CK(clk), .Q(wb_lo[5]) );
  DQV4_8TH40 wb_lo_reg_4_ ( .D(n9), .CK(clk), .Q(wb_lo[4]) );
  DQV4_8TH40 wb_lo_reg_3_ ( .D(n8), .CK(clk), .Q(wb_lo[3]) );
  DQV4_8TH40 wb_lo_reg_2_ ( .D(n7), .CK(clk), .Q(wb_lo[2]) );
  DQV4_8TH40 wb_lo_reg_1_ ( .D(n6), .CK(clk), .Q(wb_lo[1]) );
  DQV4_8TH40 wb_lo_reg_0_ ( .D(n5), .CK(clk), .Q(wb_lo[0]) );
  DQV4_8TH40 wb_hilo_we_reg ( .D(n4), .CK(clk), .Q(wb_hilo_we) );
  DQV4_8TH40 wb_llbit_we_reg ( .D(n3), .CK(clk), .Q(wb_llbit_we) );
  DQV4_8TH40 wb_llbit_value_reg ( .D(n2), .CK(clk), .Q(wb_llbit_value) );
  INOR2V4_8TH40 U2 ( .A1(mem_llbit_we), .B1(n1), .ZN(n3) );
  INOR2V0_8TH40 U3 ( .A1(mem_llbit_value), .B1(n1), .ZN(n2) );
  INOR2V0_8TH40 U4 ( .A1(mem_hilo_we), .B1(n1), .ZN(n4) );
  INOR2V0_8TH40 U5 ( .A1(mem_lo[0]), .B1(n1), .ZN(n5) );
  INOR2V0_8TH40 U6 ( .A1(mem_lo[1]), .B1(n1), .ZN(n6) );
  INOR2V0_8TH40 U7 ( .A1(mem_lo[2]), .B1(n1), .ZN(n7) );
  INOR2V0_8TH40 U8 ( .A1(mem_lo[3]), .B1(n1), .ZN(n8) );
  INOR2V0_8TH40 U9 ( .A1(mem_lo[4]), .B1(n1), .ZN(n9) );
  INOR2V0_8TH40 U10 ( .A1(mem_lo[5]), .B1(n1), .ZN(n10) );
  INOR2V0_8TH40 U11 ( .A1(mem_lo[6]), .B1(n1), .ZN(n11) );
  INOR2V0_8TH40 U12 ( .A1(mem_lo[7]), .B1(n1), .ZN(n12) );
  INOR2V0_8TH40 U13 ( .A1(mem_lo[8]), .B1(n1), .ZN(n13) );
  INOR2V0_8TH40 U14 ( .A1(mem_lo[9]), .B1(n1), .ZN(n14) );
  INOR2V0_8TH40 U15 ( .A1(mem_lo[10]), .B1(n1), .ZN(n15) );
  INOR2V0_8TH40 U16 ( .A1(mem_lo[11]), .B1(n1), .ZN(n16) );
  INOR2V0_8TH40 U17 ( .A1(mem_lo[12]), .B1(n1), .ZN(n17) );
  INOR2V0_8TH40 U18 ( .A1(mem_lo[13]), .B1(n1), .ZN(n18) );
  INOR2V0_8TH40 U19 ( .A1(mem_lo[14]), .B1(n1), .ZN(n19) );
  INOR2V0_8TH40 U20 ( .A1(mem_lo[15]), .B1(n1), .ZN(n20) );
  INOR2V0_8TH40 U21 ( .A1(mem_lo[16]), .B1(n1), .ZN(n21) );
  INOR2V0_8TH40 U22 ( .A1(mem_lo[17]), .B1(n1), .ZN(n22) );
  INOR2V0_8TH40 U23 ( .A1(mem_lo[18]), .B1(n1), .ZN(n23) );
  INOR2V0_8TH40 U24 ( .A1(mem_lo[19]), .B1(n1), .ZN(n24) );
  INOR2V0_8TH40 U25 ( .A1(mem_lo[20]), .B1(n1), .ZN(n25) );
  INOR2V0_8TH40 U26 ( .A1(mem_lo[21]), .B1(n1), .ZN(n26) );
  INOR2V0_8TH40 U27 ( .A1(mem_lo[22]), .B1(n1), .ZN(n27) );
  INOR2V0_8TH40 U28 ( .A1(mem_lo[23]), .B1(n1), .ZN(n28) );
  INOR2V0_8TH40 U29 ( .A1(mem_lo[24]), .B1(n1), .ZN(n29) );
  INOR2V0_8TH40 U30 ( .A1(mem_lo[25]), .B1(n1), .ZN(n30) );
  INOR2V0_8TH40 U31 ( .A1(mem_lo[26]), .B1(n1), .ZN(n31) );
  INOR2V0_8TH40 U32 ( .A1(mem_lo[27]), .B1(n1), .ZN(n32) );
  INOR2V0_8TH40 U33 ( .A1(mem_lo[28]), .B1(n1), .ZN(n33) );
  INOR2V0_8TH40 U34 ( .A1(mem_lo[29]), .B1(n1), .ZN(n34) );
  INOR2V0_8TH40 U35 ( .A1(mem_lo[30]), .B1(n1), .ZN(n35) );
  INOR2V0_8TH40 U36 ( .A1(mem_lo[31]), .B1(n1), .ZN(n36) );
  INOR2V0_8TH40 U37 ( .A1(mem_hi[0]), .B1(n1), .ZN(n37) );
  INOR2V0_8TH40 U38 ( .A1(mem_hi[1]), .B1(n1), .ZN(n38) );
  INOR2V0_8TH40 U39 ( .A1(mem_hi[2]), .B1(n1), .ZN(n39) );
  INOR2V0_8TH40 U40 ( .A1(mem_hi[3]), .B1(n1), .ZN(n40) );
  INOR2V0_8TH40 U41 ( .A1(mem_hi[4]), .B1(n1), .ZN(n41) );
  INOR2V0_8TH40 U42 ( .A1(mem_hi[5]), .B1(n1), .ZN(n42) );
  INOR2V0_8TH40 U43 ( .A1(mem_hi[6]), .B1(n1), .ZN(n43) );
  INOR2V0_8TH40 U44 ( .A1(mem_hi[7]), .B1(n1), .ZN(n44) );
  INOR2V0_8TH40 U45 ( .A1(mem_hi[8]), .B1(n1), .ZN(n45) );
  INOR2V0_8TH40 U46 ( .A1(mem_hi[9]), .B1(n1), .ZN(n46) );
  INOR2V0_8TH40 U47 ( .A1(mem_hi[10]), .B1(n1), .ZN(n47) );
  INOR2V0_8TH40 U48 ( .A1(mem_hi[11]), .B1(n1), .ZN(n48) );
  INOR2V0_8TH40 U49 ( .A1(mem_hi[12]), .B1(n1), .ZN(n49) );
  INOR2V0_8TH40 U50 ( .A1(mem_hi[13]), .B1(n1), .ZN(n50) );
  INOR2V0_8TH40 U51 ( .A1(mem_hi[14]), .B1(n1), .ZN(n51) );
  INOR2V0_8TH40 U52 ( .A1(mem_hi[15]), .B1(n1), .ZN(n52) );
  INOR2V0_8TH40 U53 ( .A1(mem_hi[16]), .B1(n1), .ZN(n53) );
  INOR2V0_8TH40 U54 ( .A1(mem_hi[17]), .B1(n1), .ZN(n54) );
  INOR2V0_8TH40 U55 ( .A1(mem_hi[18]), .B1(n1), .ZN(n55) );
  INOR2V0_8TH40 U56 ( .A1(mem_hi[19]), .B1(n1), .ZN(n56) );
  INOR2V0_8TH40 U57 ( .A1(mem_hi[20]), .B1(n1), .ZN(n57) );
  INOR2V0_8TH40 U58 ( .A1(mem_hi[21]), .B1(n1), .ZN(n58) );
  INOR2V0_8TH40 U59 ( .A1(mem_hi[22]), .B1(n1), .ZN(n59) );
  INOR2V0_8TH40 U60 ( .A1(mem_hi[23]), .B1(n1), .ZN(n60) );
  INOR2V0_8TH40 U61 ( .A1(mem_hi[24]), .B1(n1), .ZN(n61) );
  INOR2V0_8TH40 U62 ( .A1(mem_hi[25]), .B1(n1), .ZN(n62) );
  INOR2V0_8TH40 U63 ( .A1(mem_hi[26]), .B1(n1), .ZN(n63) );
  INOR2V0_8TH40 U64 ( .A1(mem_hi[27]), .B1(n1), .ZN(n64) );
  INOR2V0_8TH40 U65 ( .A1(mem_hi[28]), .B1(n1), .ZN(n65) );
  INOR2V0_8TH40 U66 ( .A1(mem_hi[29]), .B1(n1), .ZN(n66) );
  INOR2V0_8TH40 U67 ( .A1(mem_hi[30]), .B1(n1), .ZN(n67) );
  INOR2V0_8TH40 U68 ( .A1(mem_hi[31]), .B1(n1), .ZN(n68) );
  INOR2V0_8TH40 U69 ( .A1(mem_exe_result[0]), .B1(n1), .ZN(n69) );
  INOR2V0_8TH40 U70 ( .A1(mem_exe_result[1]), .B1(n1), .ZN(n70) );
  INOR2V0_8TH40 U71 ( .A1(mem_exe_result[2]), .B1(n1), .ZN(n71) );
  INOR2V0_8TH40 U72 ( .A1(mem_exe_result[3]), .B1(n1), .ZN(n72) );
  INOR2V0_8TH40 U73 ( .A1(mem_exe_result[4]), .B1(n1), .ZN(n73) );
  INOR2V0_8TH40 U74 ( .A1(mem_exe_result[5]), .B1(n1), .ZN(n74) );
  INOR2V0_8TH40 U75 ( .A1(mem_exe_result[6]), .B1(n1), .ZN(n75) );
  INOR2V0_8TH40 U76 ( .A1(mem_exe_result[7]), .B1(n1), .ZN(n76) );
  INOR2V0_8TH40 U77 ( .A1(mem_exe_result[8]), .B1(n1), .ZN(n77) );
  INOR2V0_8TH40 U78 ( .A1(mem_exe_result[9]), .B1(n1), .ZN(n78) );
  INOR2V0_8TH40 U79 ( .A1(mem_exe_result[10]), .B1(n1), .ZN(n79) );
  INOR2V0_8TH40 U80 ( .A1(mem_exe_result[11]), .B1(n1), .ZN(n80) );
  INOR2V0_8TH40 U81 ( .A1(mem_exe_result[12]), .B1(n1), .ZN(n81) );
  INOR2V0_8TH40 U82 ( .A1(mem_exe_result[13]), .B1(n1), .ZN(n82) );
  INOR2V0_8TH40 U83 ( .A1(mem_exe_result[14]), .B1(n1), .ZN(n83) );
  INOR2V0_8TH40 U84 ( .A1(mem_exe_result[15]), .B1(n1), .ZN(n84) );
  INOR2V0_8TH40 U85 ( .A1(mem_exe_result[16]), .B1(n1), .ZN(n85) );
  INOR2V0_8TH40 U86 ( .A1(mem_exe_result[17]), .B1(n1), .ZN(n86) );
  INOR2V0_8TH40 U87 ( .A1(mem_exe_result[18]), .B1(n1), .ZN(n87) );
  INOR2V0_8TH40 U88 ( .A1(mem_exe_result[19]), .B1(n1), .ZN(n88) );
  INOR2V0_8TH40 U89 ( .A1(mem_exe_result[20]), .B1(n1), .ZN(n89) );
  INOR2V0_8TH40 U90 ( .A1(mem_exe_result[21]), .B1(n1), .ZN(n90) );
  INOR2V0_8TH40 U91 ( .A1(mem_exe_result[22]), .B1(n1), .ZN(n91) );
  INOR2V0_8TH40 U92 ( .A1(mem_exe_result[23]), .B1(n1), .ZN(n92) );
  INOR2V0_8TH40 U93 ( .A1(mem_exe_result[24]), .B1(n1), .ZN(n93) );
  INOR2V0_8TH40 U94 ( .A1(mem_exe_result[25]), .B1(n1), .ZN(n94) );
  INOR2V0_8TH40 U95 ( .A1(mem_exe_result[26]), .B1(n1), .ZN(n95) );
  INOR2V0_8TH40 U96 ( .A1(mem_exe_result[27]), .B1(n1), .ZN(n96) );
  INOR2V0_8TH40 U97 ( .A1(mem_exe_result[28]), .B1(n1), .ZN(n97) );
  INOR2V0_8TH40 U98 ( .A1(mem_exe_result[29]), .B1(n1), .ZN(n98) );
  INOR2V0_8TH40 U99 ( .A1(mem_exe_result[30]), .B1(n1), .ZN(n99) );
  INOR2V0_8TH40 U100 ( .A1(mem_exe_result[31]), .B1(n1), .ZN(n100) );
  INOR2V0_8TH40 U101 ( .A1(mem_target_gpr[0]), .B1(n1), .ZN(n101) );
  INOR2V0_8TH40 U102 ( .A1(mem_target_gpr[1]), .B1(n1), .ZN(n102) );
  INOR2V0_8TH40 U103 ( .A1(mem_target_gpr[2]), .B1(n1), .ZN(n103) );
  INOR2V0_8TH40 U104 ( .A1(mem_target_gpr[3]), .B1(n1), .ZN(n104) );
  INOR2V0_8TH40 U105 ( .A1(mem_target_gpr[4]), .B1(n1), .ZN(n105) );
  INOR2V0_8TH40 U106 ( .A1(mem_gpr_we), .B1(n1), .ZN(n106) );
  INOR2V0_8TH40 U107 ( .A1(mem_cp0_wdata[0]), .B1(n1), .ZN(n107) );
  INOR2V0_8TH40 U108 ( .A1(mem_cp0_wdata[1]), .B1(n1), .ZN(n108) );
  INOR2V0_8TH40 U109 ( .A1(mem_cp0_wdata[2]), .B1(n1), .ZN(n109) );
  INOR2V0_8TH40 U110 ( .A1(mem_cp0_wdata[3]), .B1(n1), .ZN(n110) );
  INOR2V0_8TH40 U111 ( .A1(mem_cp0_wdata[4]), .B1(n1), .ZN(n111) );
  INOR2V0_8TH40 U112 ( .A1(mem_cp0_wdata[5]), .B1(n1), .ZN(n112) );
  INOR2V0_8TH40 U113 ( .A1(mem_cp0_wdata[6]), .B1(n1), .ZN(n113) );
  INOR2V0_8TH40 U114 ( .A1(mem_cp0_wdata[7]), .B1(n1), .ZN(n114) );
  INOR2V0_8TH40 U115 ( .A1(mem_cp0_wdata[8]), .B1(n1), .ZN(n115) );
  INOR2V0_8TH40 U116 ( .A1(mem_cp0_wdata[9]), .B1(n1), .ZN(n116) );
  INOR2V0_8TH40 U117 ( .A1(mem_cp0_wdata[10]), .B1(n1), .ZN(n117) );
  INOR2V0_8TH40 U118 ( .A1(mem_cp0_wdata[11]), .B1(n1), .ZN(n118) );
  INOR2V0_8TH40 U119 ( .A1(mem_cp0_wdata[12]), .B1(n1), .ZN(n119) );
  INOR2V0_8TH40 U120 ( .A1(mem_cp0_wdata[13]), .B1(n1), .ZN(n120) );
  INOR2V0_8TH40 U121 ( .A1(mem_cp0_wdata[14]), .B1(n1), .ZN(n121) );
  INOR2V0_8TH40 U122 ( .A1(mem_cp0_wdata[15]), .B1(n1), .ZN(n122) );
  INOR2V0_8TH40 U123 ( .A1(mem_cp0_wdata[16]), .B1(n1), .ZN(n123) );
  INOR2V0_8TH40 U124 ( .A1(mem_cp0_wdata[17]), .B1(n1), .ZN(n124) );
  INOR2V0_8TH40 U125 ( .A1(mem_cp0_wdata[18]), .B1(n1), .ZN(n125) );
  INOR2V0_8TH40 U126 ( .A1(mem_cp0_wdata[19]), .B1(n1), .ZN(n126) );
  INOR2V0_8TH40 U127 ( .A1(mem_cp0_wdata[20]), .B1(n1), .ZN(n127) );
  INOR2V0_8TH40 U128 ( .A1(mem_cp0_wdata[21]), .B1(n1), .ZN(n128) );
  INOR2V0_8TH40 U129 ( .A1(mem_cp0_wdata[22]), .B1(n1), .ZN(n129) );
  INOR2V0_8TH40 U130 ( .A1(mem_cp0_wdata[23]), .B1(n1), .ZN(n130) );
  INOR2V0_8TH40 U131 ( .A1(mem_cp0_wdata[24]), .B1(n1), .ZN(n131) );
  INOR2V0_8TH40 U132 ( .A1(mem_cp0_wdata[25]), .B1(n1), .ZN(n132) );
  INOR2V0_8TH40 U133 ( .A1(mem_cp0_wdata[26]), .B1(n1), .ZN(n133) );
  INOR2V0_8TH40 U134 ( .A1(mem_cp0_wdata[27]), .B1(n1), .ZN(n134) );
  INOR2V0_8TH40 U135 ( .A1(mem_cp0_wdata[28]), .B1(n1), .ZN(n135) );
  INOR2V0_8TH40 U136 ( .A1(mem_cp0_wdata[29]), .B1(n1), .ZN(n136) );
  INOR2V0_8TH40 U137 ( .A1(mem_cp0_wdata[30]), .B1(n1), .ZN(n137) );
  INOR2V0_8TH40 U138 ( .A1(mem_cp0_wdata[31]), .B1(n1), .ZN(n138) );
  INOR2V0_8TH40 U139 ( .A1(mem_cp0_waddr[0]), .B1(n1), .ZN(n139) );
  INOR2V0_8TH40 U140 ( .A1(mem_cp0_waddr[1]), .B1(n1), .ZN(n140) );
  INOR2V0_8TH40 U141 ( .A1(mem_cp0_waddr[2]), .B1(n1), .ZN(n141) );
  INOR2V0_8TH40 U142 ( .A1(mem_cp0_waddr[3]), .B1(n1), .ZN(n142) );
  INOR2V0_8TH40 U143 ( .A1(mem_cp0_waddr[4]), .B1(n1), .ZN(n143) );
  INOR2V0_8TH40 U144 ( .A1(mem_cp0_we), .B1(n1), .ZN(n144) );
  I2NAND3V1_8TH40 U145 ( .A1(stall_ctrl[4]), .A2(rst), .B(flush_BAR), .ZN(n1)
         );
endmodule


module hilo_reg ( clk, rst, we, hi_i, lo_i, hi_o, lo_o );
  input [31:0] hi_i;
  input [31:0] lo_i;
  output [31:0] hi_o;
  output [31:0] lo_o;
  input clk, rst, we;
  wire   n1;

  EDGRNQV2_8TH40 lo_o_reg_31_ ( .RN(n1), .D(lo_i[31]), .E(we), .CK(clk), .Q(
        lo_o[31]) );
  EDGRNQV2_8TH40 lo_o_reg_29_ ( .RN(n1), .D(lo_i[29]), .E(we), .CK(clk), .Q(
        lo_o[29]) );
  EDGRNQV2_8TH40 lo_o_reg_27_ ( .RN(n1), .D(lo_i[27]), .E(we), .CK(clk), .Q(
        lo_o[27]) );
  EDGRNQV2_8TH40 lo_o_reg_26_ ( .RN(n1), .D(lo_i[26]), .E(we), .CK(clk), .Q(
        lo_o[26]) );
  EDGRNQV2_8TH40 lo_o_reg_25_ ( .RN(n1), .D(lo_i[25]), .E(we), .CK(clk), .Q(
        lo_o[25]) );
  EDGRNQV2_8TH40 lo_o_reg_24_ ( .RN(n1), .D(lo_i[24]), .E(we), .CK(clk), .Q(
        lo_o[24]) );
  EDGRNQV2_8TH40 lo_o_reg_23_ ( .RN(n1), .D(lo_i[23]), .E(we), .CK(clk), .Q(
        lo_o[23]) );
  EDGRNQV2_8TH40 lo_o_reg_22_ ( .RN(n1), .D(lo_i[22]), .E(we), .CK(clk), .Q(
        lo_o[22]) );
  EDGRNQV2_8TH40 lo_o_reg_20_ ( .RN(n1), .D(lo_i[20]), .E(we), .CK(clk), .Q(
        lo_o[20]) );
  EDGRNQV2_8TH40 lo_o_reg_19_ ( .RN(n1), .D(lo_i[19]), .E(we), .CK(clk), .Q(
        lo_o[19]) );
  EDGRNQV2_8TH40 lo_o_reg_15_ ( .RN(n1), .D(lo_i[15]), .E(we), .CK(clk), .Q(
        lo_o[15]) );
  EDGRNQV2_8TH40 lo_o_reg_14_ ( .RN(n1), .D(lo_i[14]), .E(we), .CK(clk), .Q(
        lo_o[14]) );
  EDGRNQV2_8TH40 lo_o_reg_12_ ( .RN(n1), .D(lo_i[12]), .E(we), .CK(clk), .Q(
        lo_o[12]) );
  EDGRNQV2_8TH40 lo_o_reg_7_ ( .RN(n1), .D(lo_i[7]), .E(we), .CK(clk), .Q(
        lo_o[7]) );
  EDGRNQV2_8TH40 lo_o_reg_5_ ( .RN(n1), .D(lo_i[5]), .E(we), .CK(clk), .Q(
        lo_o[5]) );
  EDGRNQV2_8TH40 lo_o_reg_3_ ( .RN(n1), .D(lo_i[3]), .E(we), .CK(clk), .Q(
        lo_o[3]) );
  EDGRNQV2_8TH40 lo_o_reg_0_ ( .RN(n1), .D(lo_i[0]), .E(we), .CK(clk), .Q(
        lo_o[0]) );
  EDGRNQV2_8TH40 lo_o_reg_30_ ( .RN(n1), .D(lo_i[30]), .E(we), .CK(clk), .Q(
        lo_o[30]) );
  EDGRNQV2_8TH40 lo_o_reg_28_ ( .RN(n1), .D(lo_i[28]), .E(we), .CK(clk), .Q(
        lo_o[28]) );
  EDGRNQV2_8TH40 lo_o_reg_21_ ( .RN(n1), .D(lo_i[21]), .E(we), .CK(clk), .Q(
        lo_o[21]) );
  EDGRNQV2_8TH40 lo_o_reg_18_ ( .RN(n1), .D(lo_i[18]), .E(we), .CK(clk), .Q(
        lo_o[18]) );
  EDGRNQV2_8TH40 lo_o_reg_17_ ( .RN(n1), .D(lo_i[17]), .E(we), .CK(clk), .Q(
        lo_o[17]) );
  EDGRNQV2_8TH40 lo_o_reg_16_ ( .RN(n1), .D(lo_i[16]), .E(we), .CK(clk), .Q(
        lo_o[16]) );
  EDGRNQV2_8TH40 lo_o_reg_13_ ( .RN(n1), .D(lo_i[13]), .E(we), .CK(clk), .Q(
        lo_o[13]) );
  EDGRNQV2_8TH40 lo_o_reg_11_ ( .RN(n1), .D(lo_i[11]), .E(we), .CK(clk), .Q(
        lo_o[11]) );
  EDGRNQV2_8TH40 lo_o_reg_10_ ( .RN(n1), .D(lo_i[10]), .E(we), .CK(clk), .Q(
        lo_o[10]) );
  EDGRNQV2_8TH40 lo_o_reg_9_ ( .RN(n1), .D(lo_i[9]), .E(we), .CK(clk), .Q(
        lo_o[9]) );
  EDGRNQV2_8TH40 lo_o_reg_8_ ( .RN(n1), .D(lo_i[8]), .E(we), .CK(clk), .Q(
        lo_o[8]) );
  EDGRNQV2_8TH40 lo_o_reg_6_ ( .RN(n1), .D(lo_i[6]), .E(we), .CK(clk), .Q(
        lo_o[6]) );
  EDGRNQV2_8TH40 lo_o_reg_4_ ( .RN(n1), .D(lo_i[4]), .E(we), .CK(clk), .Q(
        lo_o[4]) );
  EDGRNQV2_8TH40 lo_o_reg_2_ ( .RN(n1), .D(lo_i[2]), .E(we), .CK(clk), .Q(
        lo_o[2]) );
  EDGRNQV2_8TH40 lo_o_reg_1_ ( .RN(n1), .D(lo_i[1]), .E(we), .CK(clk), .Q(
        lo_o[1]) );
  EDGRNQV2_8TH40 hi_o_reg_31_ ( .RN(n1), .D(hi_i[31]), .E(we), .CK(clk), .Q(
        hi_o[31]) );
  EDGRNQV2_8TH40 hi_o_reg_30_ ( .RN(n1), .D(hi_i[30]), .E(we), .CK(clk), .Q(
        hi_o[30]) );
  EDGRNQV2_8TH40 hi_o_reg_29_ ( .RN(n1), .D(hi_i[29]), .E(we), .CK(clk), .Q(
        hi_o[29]) );
  EDGRNQV2_8TH40 hi_o_reg_28_ ( .RN(n1), .D(hi_i[28]), .E(we), .CK(clk), .Q(
        hi_o[28]) );
  EDGRNQV2_8TH40 hi_o_reg_27_ ( .RN(n1), .D(hi_i[27]), .E(we), .CK(clk), .Q(
        hi_o[27]) );
  EDGRNQV2_8TH40 hi_o_reg_26_ ( .RN(n1), .D(hi_i[26]), .E(we), .CK(clk), .Q(
        hi_o[26]) );
  EDGRNQV2_8TH40 hi_o_reg_25_ ( .RN(n1), .D(hi_i[25]), .E(we), .CK(clk), .Q(
        hi_o[25]) );
  EDGRNQV2_8TH40 hi_o_reg_24_ ( .RN(n1), .D(hi_i[24]), .E(we), .CK(clk), .Q(
        hi_o[24]) );
  EDGRNQV2_8TH40 hi_o_reg_23_ ( .RN(n1), .D(hi_i[23]), .E(we), .CK(clk), .Q(
        hi_o[23]) );
  EDGRNQV2_8TH40 hi_o_reg_22_ ( .RN(n1), .D(hi_i[22]), .E(we), .CK(clk), .Q(
        hi_o[22]) );
  EDGRNQV2_8TH40 hi_o_reg_21_ ( .RN(n1), .D(hi_i[21]), .E(we), .CK(clk), .Q(
        hi_o[21]) );
  EDGRNQV2_8TH40 hi_o_reg_20_ ( .RN(n1), .D(hi_i[20]), .E(we), .CK(clk), .Q(
        hi_o[20]) );
  EDGRNQV2_8TH40 hi_o_reg_19_ ( .RN(n1), .D(hi_i[19]), .E(we), .CK(clk), .Q(
        hi_o[19]) );
  EDGRNQV2_8TH40 hi_o_reg_18_ ( .RN(n1), .D(hi_i[18]), .E(we), .CK(clk), .Q(
        hi_o[18]) );
  EDGRNQV2_8TH40 hi_o_reg_17_ ( .RN(n1), .D(hi_i[17]), .E(we), .CK(clk), .Q(
        hi_o[17]) );
  EDGRNQV2_8TH40 hi_o_reg_16_ ( .RN(n1), .D(hi_i[16]), .E(we), .CK(clk), .Q(
        hi_o[16]) );
  EDGRNQV2_8TH40 hi_o_reg_15_ ( .RN(n1), .D(hi_i[15]), .E(we), .CK(clk), .Q(
        hi_o[15]) );
  EDGRNQV2_8TH40 hi_o_reg_14_ ( .RN(n1), .D(hi_i[14]), .E(we), .CK(clk), .Q(
        hi_o[14]) );
  EDGRNQV2_8TH40 hi_o_reg_13_ ( .RN(n1), .D(hi_i[13]), .E(we), .CK(clk), .Q(
        hi_o[13]) );
  EDGRNQV2_8TH40 hi_o_reg_12_ ( .RN(n1), .D(hi_i[12]), .E(we), .CK(clk), .Q(
        hi_o[12]) );
  EDGRNQV2_8TH40 hi_o_reg_11_ ( .RN(n1), .D(hi_i[11]), .E(we), .CK(clk), .Q(
        hi_o[11]) );
  EDGRNQV2_8TH40 hi_o_reg_10_ ( .RN(n1), .D(hi_i[10]), .E(we), .CK(clk), .Q(
        hi_o[10]) );
  EDGRNQV2_8TH40 hi_o_reg_9_ ( .RN(n1), .D(hi_i[9]), .E(we), .CK(clk), .Q(
        hi_o[9]) );
  EDGRNQV2_8TH40 hi_o_reg_8_ ( .RN(n1), .D(hi_i[8]), .E(we), .CK(clk), .Q(
        hi_o[8]) );
  EDGRNQV2_8TH40 hi_o_reg_7_ ( .RN(n1), .D(hi_i[7]), .E(we), .CK(clk), .Q(
        hi_o[7]) );
  EDGRNQV2_8TH40 hi_o_reg_6_ ( .RN(n1), .D(hi_i[6]), .E(we), .CK(clk), .Q(
        hi_o[6]) );
  EDGRNQV2_8TH40 hi_o_reg_5_ ( .RN(n1), .D(hi_i[5]), .E(we), .CK(clk), .Q(
        hi_o[5]) );
  EDGRNQV2_8TH40 hi_o_reg_4_ ( .RN(n1), .D(hi_i[4]), .E(we), .CK(clk), .Q(
        hi_o[4]) );
  EDGRNQV2_8TH40 hi_o_reg_3_ ( .RN(n1), .D(hi_i[3]), .E(we), .CK(clk), .Q(
        hi_o[3]) );
  EDGRNQV2_8TH40 hi_o_reg_2_ ( .RN(n1), .D(hi_i[2]), .E(we), .CK(clk), .Q(
        hi_o[2]) );
  EDGRNQV2_8TH40 hi_o_reg_1_ ( .RN(n1), .D(hi_i[1]), .E(we), .CK(clk), .Q(
        hi_o[1]) );
  EDGRNQV2_8TH40 hi_o_reg_0_ ( .RN(n1), .D(hi_i[0]), .E(we), .CK(clk), .Q(
        hi_o[0]) );
  CLKNV1_8TH40 U2 ( .I(rst), .ZN(n1) );
endmodule


module llbit_reg ( clk, rst, we, llbit_i, llbit_o, flush_BAR );
  input clk, rst, we, llbit_i, flush_BAR;
  output llbit_o;
  wire   n3, n1;

  DQV4_8TH40 llbit_o_reg ( .D(n3), .CK(clk), .Q(llbit_o) );
  INOR3V2_8TH40 U2 ( .A1(flush_BAR), .B1(n1), .B2(rst), .ZN(n3) );
  MUX2NV0_8TH40 U3 ( .I0(llbit_o), .I1(llbit_i), .S(we), .ZN(n1) );
endmodule


module pipe_ctrl ( rst, stall_req_if, stall_req_id, stall_req_ex, 
        stall_req_mem, cp0_epc, except_type, pc_new, stall_ctrl, flush_BAR );
  input [31:0] cp0_epc;
  input [31:0] except_type;
  output [31:0] pc_new;
  output [5:0] stall_ctrl;
  input rst, stall_req_if, stall_req_id, stall_req_ex, stall_req_mem;
  output flush_BAR;
  wire   N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  assign stall_ctrl[0] = stall_ctrl[2];
  assign stall_ctrl[1] = stall_ctrl[2];

  LAHQV1_8TH40 pc_new_reg_3_ ( .E(N124), .D(N128), .Q(pc_new[3]) );
  LAHQV1_8TH40 pc_new_reg_2_ ( .E(N124), .D(N127), .Q(pc_new[2]) );
  LAHQV1_8TH40 pc_new_reg_1_ ( .E(N124), .D(N126), .Q(pc_new[1]) );
  LAHQV1_8TH40 pc_new_reg_0_ ( .E(N124), .D(N125), .Q(pc_new[0]) );
  LAHQV4_8TH40 pc_new_reg_31_ ( .E(N124), .D(N156), .Q(pc_new[31]) );
  LAHQV4_8TH40 pc_new_reg_30_ ( .E(N124), .D(N155), .Q(pc_new[30]) );
  LAHQV4_8TH40 pc_new_reg_29_ ( .E(N124), .D(N154), .Q(pc_new[29]) );
  LAHQV4_8TH40 pc_new_reg_28_ ( .E(N124), .D(N153), .Q(pc_new[28]) );
  LAHQV4_8TH40 pc_new_reg_27_ ( .E(N124), .D(N152), .Q(pc_new[27]) );
  LAHQV4_8TH40 pc_new_reg_26_ ( .E(N124), .D(N151), .Q(pc_new[26]) );
  LAHQV4_8TH40 pc_new_reg_25_ ( .E(N124), .D(N150), .Q(pc_new[25]) );
  LAHQV4_8TH40 pc_new_reg_24_ ( .E(N124), .D(N149), .Q(pc_new[24]) );
  LAHQV4_8TH40 pc_new_reg_23_ ( .E(N124), .D(N148), .Q(pc_new[23]) );
  LAHQV4_8TH40 pc_new_reg_22_ ( .E(N124), .D(N147), .Q(pc_new[22]) );
  LAHQV4_8TH40 pc_new_reg_21_ ( .E(N124), .D(N146), .Q(pc_new[21]) );
  LAHQV4_8TH40 pc_new_reg_20_ ( .E(N124), .D(N145), .Q(pc_new[20]) );
  LAHQV4_8TH40 pc_new_reg_19_ ( .E(N124), .D(N144), .Q(pc_new[19]) );
  LAHQV4_8TH40 pc_new_reg_18_ ( .E(N124), .D(N143), .Q(pc_new[18]) );
  LAHQV4_8TH40 pc_new_reg_17_ ( .E(N124), .D(N142), .Q(pc_new[17]) );
  LAHQV4_8TH40 pc_new_reg_16_ ( .E(N124), .D(N141), .Q(pc_new[16]) );
  LAHQV4_8TH40 pc_new_reg_15_ ( .E(N124), .D(N140), .Q(pc_new[15]) );
  LAHQV4_8TH40 pc_new_reg_14_ ( .E(N124), .D(N139), .Q(pc_new[14]) );
  LAHQV4_8TH40 pc_new_reg_13_ ( .E(N124), .D(N138), .Q(pc_new[13]) );
  LAHQV4_8TH40 pc_new_reg_12_ ( .E(N124), .D(N137), .Q(pc_new[12]) );
  LAHQV4_8TH40 pc_new_reg_11_ ( .E(N124), .D(N136), .Q(pc_new[11]) );
  LAHQV4_8TH40 pc_new_reg_10_ ( .E(N124), .D(N135), .Q(pc_new[10]) );
  LAHQV4_8TH40 pc_new_reg_9_ ( .E(N124), .D(N134), .Q(pc_new[9]) );
  LAHQV4_8TH40 pc_new_reg_8_ ( .E(N124), .D(N133), .Q(pc_new[8]) );
  LAHQV4_8TH40 pc_new_reg_7_ ( .E(N124), .D(N132), .Q(pc_new[7]) );
  LAHQV4_8TH40 pc_new_reg_6_ ( .E(N124), .D(N131), .Q(pc_new[6]) );
  LAHQV4_8TH40 pc_new_reg_5_ ( .E(N124), .D(N130), .Q(pc_new[5]) );
  LAHQV4_8TH40 pc_new_reg_4_ ( .E(N124), .D(N129), .Q(pc_new[4]) );
  MOAI22V4_8TH40 U3 ( .A1(flush_BAR), .A2(n6), .B1(cp0_epc[5]), .B2(n4), .ZN(
        N130) );
  IOA21V8_8TH40 U4 ( .A1(cp0_epc[6]), .A2(n4), .B(n5), .ZN(N131) );
  AND2V4_8TH40 U5 ( .A1(cp0_epc[31]), .A2(n4), .Z(N156) );
  AND2V4_8TH40 U6 ( .A1(cp0_epc[30]), .A2(n4), .Z(N155) );
  AND2V4_8TH40 U7 ( .A1(cp0_epc[29]), .A2(n4), .Z(N154) );
  AND2V4_8TH40 U8 ( .A1(cp0_epc[28]), .A2(n4), .Z(N153) );
  AND2V4_8TH40 U9 ( .A1(cp0_epc[27]), .A2(n4), .Z(N152) );
  AND2V4_8TH40 U10 ( .A1(cp0_epc[26]), .A2(n4), .Z(N151) );
  AND2V4_8TH40 U11 ( .A1(cp0_epc[25]), .A2(n4), .Z(N150) );
  AND2V4_8TH40 U12 ( .A1(cp0_epc[24]), .A2(n4), .Z(N149) );
  AND2V4_8TH40 U13 ( .A1(cp0_epc[23]), .A2(n4), .Z(N148) );
  AND2V4_8TH40 U14 ( .A1(cp0_epc[22]), .A2(n4), .Z(N147) );
  AND2V4_8TH40 U15 ( .A1(cp0_epc[21]), .A2(n4), .Z(N146) );
  AND2V4_8TH40 U16 ( .A1(cp0_epc[20]), .A2(n4), .Z(N145) );
  AND2V4_8TH40 U17 ( .A1(cp0_epc[19]), .A2(n4), .Z(N144) );
  AND2V4_8TH40 U18 ( .A1(cp0_epc[18]), .A2(n4), .Z(N143) );
  AND2V4_8TH40 U19 ( .A1(cp0_epc[17]), .A2(n4), .Z(N142) );
  AND2V4_8TH40 U20 ( .A1(cp0_epc[16]), .A2(n4), .Z(N141) );
  AND2V4_8TH40 U21 ( .A1(cp0_epc[15]), .A2(n4), .Z(N140) );
  AND2V4_8TH40 U22 ( .A1(cp0_epc[14]), .A2(n4), .Z(N139) );
  AND2V4_8TH40 U23 ( .A1(cp0_epc[13]), .A2(n4), .Z(N138) );
  AND2V4_8TH40 U24 ( .A1(cp0_epc[12]), .A2(n4), .Z(N137) );
  AND2V4_8TH40 U25 ( .A1(cp0_epc[11]), .A2(n4), .Z(N136) );
  AND2V4_8TH40 U26 ( .A1(cp0_epc[10]), .A2(n4), .Z(N135) );
  AND2V4_8TH40 U27 ( .A1(cp0_epc[9]), .A2(n4), .Z(N134) );
  AND2V4_8TH40 U28 ( .A1(cp0_epc[8]), .A2(n4), .Z(N133) );
  AND2V4_8TH40 U29 ( .A1(cp0_epc[7]), .A2(n4), .Z(N132) );
  AND2V4_8TH40 U30 ( .A1(cp0_epc[4]), .A2(n4), .Z(N129) );
  AND2V4_8TH40 U31 ( .A1(cp0_epc[3]), .A2(n4), .Z(N128) );
  AND2V4_8TH40 U32 ( .A1(cp0_epc[2]), .A2(n4), .Z(N127) );
  AND2V4_8TH40 U33 ( .A1(cp0_epc[1]), .A2(n4), .Z(N126) );
  AND2V4_8TH40 U34 ( .A1(cp0_epc[0]), .A2(n4), .Z(N125) );
  NAND3V2_8TH40 U35 ( .A1(except_type[3]), .A2(n8), .A3(n12), .ZN(n5) );
  I2NAND4V2_8TH40 U36 ( .A1(flush_BAR), .A2(except_type[0]), .B1(n9), .B2(
        except_type[1]), .ZN(n7) );
  OAO211V2_8TH40 U37 ( .A1(stall_req_id), .A2(stall_req_if), .B(n2), .C(
        stall_ctrl[3]), .Z(stall_ctrl[2]) );
  NAND2V2_8TH40 U38 ( .A1(stall_req_mem), .A2(n2), .ZN(n1) );
  CLKNV1_8TH40 U39 ( .I(n1), .ZN(stall_ctrl[4]) );
  IOA21V0_8TH40 U40 ( .A1(stall_req_ex), .A2(n2), .B(n1), .ZN(stall_ctrl[3])
         );
  INOR2V0_8TH40 U41 ( .A1(n3), .B1(rst), .ZN(n2) );
  CLKNV1_8TH40 U42 ( .I(n7), .ZN(n4) );
  NAND4V0P5_8TH40 U43 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(N124) );
  NOR2V0P5_8TH40 U44 ( .A1(n10), .A2(n11), .ZN(n9) );
  CLKNV1_8TH40 U45 ( .I(n8), .ZN(flush_BAR) );
  I2NAND3V1_8TH40 U46 ( .A1(except_type[1]), .A2(except_type[2]), .B(n11), 
        .ZN(n6) );
  CLKNV1_8TH40 U47 ( .I(except_type[3]), .ZN(n11) );
  MUX2NV0_8TH40 U48 ( .I0(except_type[1]), .I1(except_type[0]), .S(n10), .ZN(
        n12) );
  CLKNV1_8TH40 U49 ( .I(except_type[2]), .ZN(n10) );
  NOR2V0P5_8TH40 U50 ( .A1(rst), .A2(n3), .ZN(n8) );
  NOR4V0P5_8TH40 U51 ( .A1(except_type[0]), .A2(except_type[1]), .A3(
        except_type[2]), .A4(except_type[3]), .ZN(n3) );
endmodule


module div_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62;
  assign DIFF[0] = B[0];

  AND2V2_8TH40 U1 ( .A1(n31), .A2(n42), .Z(n1) );
  AND2V2_8TH40 U2 ( .A1(n1), .A2(n53), .Z(n2) );
  AND2V2_8TH40 U3 ( .A1(n2), .A2(n56), .Z(n3) );
  AND2V2_8TH40 U4 ( .A1(n3), .A2(n57), .Z(n4) );
  AND2V2_8TH40 U5 ( .A1(n4), .A2(n58), .Z(n5) );
  AND2V2_8TH40 U6 ( .A1(n5), .A2(n59), .Z(n6) );
  AND2V2_8TH40 U7 ( .A1(n6), .A2(n60), .Z(n7) );
  AND2V2_8TH40 U8 ( .A1(n7), .A2(n61), .Z(n8) );
  AND2V2_8TH40 U9 ( .A1(n8), .A2(n62), .Z(n9) );
  AND2V2_8TH40 U10 ( .A1(n9), .A2(n32), .Z(n10) );
  AND2V2_8TH40 U11 ( .A1(n10), .A2(n33), .Z(n11) );
  AND2V2_8TH40 U12 ( .A1(n11), .A2(n34), .Z(n12) );
  AND2V2_8TH40 U13 ( .A1(n12), .A2(n35), .Z(n13) );
  AND2V2_8TH40 U14 ( .A1(n13), .A2(n36), .Z(n14) );
  AND2V2_8TH40 U15 ( .A1(n14), .A2(n37), .Z(n15) );
  AND2V2_8TH40 U16 ( .A1(n15), .A2(n38), .Z(n16) );
  AND2V2_8TH40 U17 ( .A1(n16), .A2(n39), .Z(n17) );
  AND2V2_8TH40 U18 ( .A1(n17), .A2(n40), .Z(n18) );
  AND2V2_8TH40 U19 ( .A1(n18), .A2(n41), .Z(n19) );
  AND2V2_8TH40 U20 ( .A1(n19), .A2(n43), .Z(n20) );
  AND2V2_8TH40 U21 ( .A1(n20), .A2(n44), .Z(n21) );
  AND2V2_8TH40 U22 ( .A1(n21), .A2(n45), .Z(n22) );
  AND2V2_8TH40 U23 ( .A1(n22), .A2(n46), .Z(n23) );
  AND2V2_8TH40 U24 ( .A1(n23), .A2(n47), .Z(n24) );
  AND2V2_8TH40 U25 ( .A1(n24), .A2(n48), .Z(n25) );
  AND2V2_8TH40 U26 ( .A1(n25), .A2(n49), .Z(n26) );
  AND2V2_8TH40 U27 ( .A1(n26), .A2(n50), .Z(n27) );
  AND2V2_8TH40 U28 ( .A1(n27), .A2(n51), .Z(n28) );
  AND2V2_8TH40 U29 ( .A1(n28), .A2(n52), .Z(n29) );
  AND2V2_8TH40 U30 ( .A1(n29), .A2(n54), .Z(n30) );
  INV2_8TH40 U31 ( .I(B[0]), .ZN(n31) );
  INV2_8TH40 U32 ( .I(B[31]), .ZN(n55) );
  INV2_8TH40 U33 ( .I(B[1]), .ZN(n42) );
  INV2_8TH40 U34 ( .I(B[2]), .ZN(n53) );
  INV2_8TH40 U35 ( .I(B[3]), .ZN(n56) );
  INV2_8TH40 U36 ( .I(B[4]), .ZN(n57) );
  INV2_8TH40 U37 ( .I(B[5]), .ZN(n58) );
  INV2_8TH40 U38 ( .I(B[6]), .ZN(n59) );
  INV2_8TH40 U39 ( .I(B[7]), .ZN(n60) );
  INV2_8TH40 U40 ( .I(B[8]), .ZN(n61) );
  INV2_8TH40 U41 ( .I(B[9]), .ZN(n62) );
  INV2_8TH40 U42 ( .I(B[10]), .ZN(n32) );
  INV2_8TH40 U43 ( .I(B[11]), .ZN(n33) );
  INV2_8TH40 U44 ( .I(B[12]), .ZN(n34) );
  INV2_8TH40 U45 ( .I(B[13]), .ZN(n35) );
  INV2_8TH40 U46 ( .I(B[14]), .ZN(n36) );
  INV2_8TH40 U47 ( .I(B[15]), .ZN(n37) );
  INV2_8TH40 U48 ( .I(B[16]), .ZN(n38) );
  INV2_8TH40 U49 ( .I(B[17]), .ZN(n39) );
  INV2_8TH40 U50 ( .I(B[18]), .ZN(n40) );
  INV2_8TH40 U51 ( .I(B[19]), .ZN(n41) );
  INV2_8TH40 U52 ( .I(B[20]), .ZN(n43) );
  INV2_8TH40 U53 ( .I(B[21]), .ZN(n44) );
  INV2_8TH40 U54 ( .I(B[22]), .ZN(n45) );
  INV2_8TH40 U55 ( .I(B[23]), .ZN(n46) );
  INV2_8TH40 U56 ( .I(B[24]), .ZN(n47) );
  INV2_8TH40 U57 ( .I(B[25]), .ZN(n48) );
  INV2_8TH40 U58 ( .I(B[26]), .ZN(n49) );
  INV2_8TH40 U59 ( .I(B[27]), .ZN(n50) );
  INV2_8TH40 U60 ( .I(B[28]), .ZN(n51) );
  INV2_8TH40 U61 ( .I(B[29]), .ZN(n52) );
  INV2_8TH40 U62 ( .I(B[30]), .ZN(n54) );
  XOR2V2_8TH40 U63 ( .A1(n55), .A2(n30), .Z(DIFF[31]) );
  XOR2V2_8TH40 U64 ( .A1(n29), .A2(n54), .Z(DIFF[30]) );
  XOR2V2_8TH40 U65 ( .A1(n28), .A2(n52), .Z(DIFF[29]) );
  XOR2V2_8TH40 U66 ( .A1(n27), .A2(n51), .Z(DIFF[28]) );
  XOR2V2_8TH40 U67 ( .A1(n26), .A2(n50), .Z(DIFF[27]) );
  XOR2V2_8TH40 U68 ( .A1(n25), .A2(n49), .Z(DIFF[26]) );
  XOR2V2_8TH40 U69 ( .A1(n24), .A2(n48), .Z(DIFF[25]) );
  XOR2V2_8TH40 U70 ( .A1(n23), .A2(n47), .Z(DIFF[24]) );
  XOR2V2_8TH40 U71 ( .A1(n22), .A2(n46), .Z(DIFF[23]) );
  XOR2V2_8TH40 U72 ( .A1(n21), .A2(n45), .Z(DIFF[22]) );
  XOR2V2_8TH40 U73 ( .A1(n20), .A2(n44), .Z(DIFF[21]) );
  XOR2V2_8TH40 U74 ( .A1(n19), .A2(n43), .Z(DIFF[20]) );
  XOR2V2_8TH40 U75 ( .A1(n18), .A2(n41), .Z(DIFF[19]) );
  XOR2V2_8TH40 U76 ( .A1(n17), .A2(n40), .Z(DIFF[18]) );
  XOR2V2_8TH40 U77 ( .A1(n16), .A2(n39), .Z(DIFF[17]) );
  XOR2V2_8TH40 U78 ( .A1(n15), .A2(n38), .Z(DIFF[16]) );
  XOR2V2_8TH40 U79 ( .A1(n14), .A2(n37), .Z(DIFF[15]) );
  XOR2V2_8TH40 U80 ( .A1(n13), .A2(n36), .Z(DIFF[14]) );
  XOR2V2_8TH40 U81 ( .A1(n12), .A2(n35), .Z(DIFF[13]) );
  XOR2V2_8TH40 U82 ( .A1(n11), .A2(n34), .Z(DIFF[12]) );
  XOR2V2_8TH40 U83 ( .A1(n10), .A2(n33), .Z(DIFF[11]) );
  XOR2V2_8TH40 U84 ( .A1(n9), .A2(n32), .Z(DIFF[10]) );
  XOR2V2_8TH40 U85 ( .A1(n8), .A2(n62), .Z(DIFF[9]) );
  XOR2V2_8TH40 U86 ( .A1(n7), .A2(n61), .Z(DIFF[8]) );
  XOR2V2_8TH40 U87 ( .A1(n6), .A2(n60), .Z(DIFF[7]) );
  XOR2V2_8TH40 U88 ( .A1(n5), .A2(n59), .Z(DIFF[6]) );
  XOR2V2_8TH40 U89 ( .A1(n4), .A2(n58), .Z(DIFF[5]) );
  XOR2V2_8TH40 U90 ( .A1(n3), .A2(n57), .Z(DIFF[4]) );
  XOR2V2_8TH40 U91 ( .A1(n2), .A2(n56), .Z(DIFF[3]) );
  XOR2V2_8TH40 U92 ( .A1(n1), .A2(n53), .Z(DIFF[2]) );
  XOR2V2_8TH40 U93 ( .A1(n31), .A2(n42), .Z(DIFF[1]) );
endmodule


module div_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;
  assign DIFF[0] = B[0];

  XOR2V4_8TH40 U1 ( .A1(B[31]), .A2(n30), .Z(DIFF[31]) );
  NAND2V2_8TH40 U2 ( .A1(n23), .A2(n54), .ZN(n30) );
  AND2V2_8TH40 U3 ( .A1(n31), .A2(n42), .Z(n1) );
  AND2V2_8TH40 U4 ( .A1(n1), .A2(n53), .Z(n2) );
  AND2V2_8TH40 U5 ( .A1(n16), .A2(n56), .Z(n3) );
  AND2V2_8TH40 U6 ( .A1(n3), .A2(n57), .Z(n4) );
  AND2V2_8TH40 U7 ( .A1(n17), .A2(n60), .Z(n5) );
  AND2V2_8TH40 U8 ( .A1(n5), .A2(n61), .Z(n6) );
  AND2V2_8TH40 U9 ( .A1(n18), .A2(n33), .Z(n7) );
  AND2V2_8TH40 U10 ( .A1(n7), .A2(n34), .Z(n8) );
  AND2V2_8TH40 U11 ( .A1(n19), .A2(n37), .Z(n9) );
  AND2V2_8TH40 U12 ( .A1(n9), .A2(n38), .Z(n10) );
  AND2V2_8TH40 U13 ( .A1(n20), .A2(n41), .Z(n11) );
  AND2V2_8TH40 U14 ( .A1(n21), .A2(n45), .Z(n12) );
  AND2V2_8TH40 U15 ( .A1(n12), .A2(n46), .Z(n13) );
  AND2V2_8TH40 U16 ( .A1(n22), .A2(n49), .Z(n14) );
  AND2V2_8TH40 U17 ( .A1(n14), .A2(n50), .Z(n15) );
  AND2V2_8TH40 U18 ( .A1(n2), .A2(n55), .Z(n16) );
  AND2V2_8TH40 U19 ( .A1(n24), .A2(n59), .Z(n17) );
  AND2V2_8TH40 U20 ( .A1(n6), .A2(n32), .Z(n18) );
  AND2V2_8TH40 U21 ( .A1(n25), .A2(n36), .Z(n19) );
  AND2V2_8TH40 U22 ( .A1(n26), .A2(n40), .Z(n20) );
  AND2V2_8TH40 U23 ( .A1(n27), .A2(n44), .Z(n21) );
  AND2V2_8TH40 U24 ( .A1(n28), .A2(n48), .Z(n22) );
  AND2V2_8TH40 U25 ( .A1(n29), .A2(n52), .Z(n23) );
  AND2V2_8TH40 U26 ( .A1(n4), .A2(n58), .Z(n24) );
  AND2V2_8TH40 U27 ( .A1(n8), .A2(n35), .Z(n25) );
  AND2V2_8TH40 U28 ( .A1(n10), .A2(n39), .Z(n26) );
  AND2V2_8TH40 U29 ( .A1(n11), .A2(n43), .Z(n27) );
  AND2V2_8TH40 U30 ( .A1(n13), .A2(n47), .Z(n28) );
  AND2V2_8TH40 U31 ( .A1(n15), .A2(n51), .Z(n29) );
  INV2_8TH40 U32 ( .I(B[0]), .ZN(n31) );
  INV2_8TH40 U33 ( .I(B[2]), .ZN(n53) );
  INV2_8TH40 U34 ( .I(B[4]), .ZN(n56) );
  INV2_8TH40 U35 ( .I(B[8]), .ZN(n60) );
  INV2_8TH40 U36 ( .I(B[11]), .ZN(n33) );
  INV2_8TH40 U37 ( .I(B[15]), .ZN(n37) );
  INV2_8TH40 U38 ( .I(B[19]), .ZN(n41) );
  INV2_8TH40 U39 ( .I(B[22]), .ZN(n45) );
  INV2_8TH40 U40 ( .I(B[26]), .ZN(n49) );
  INV2_8TH40 U41 ( .I(B[1]), .ZN(n42) );
  INV2_8TH40 U42 ( .I(B[5]), .ZN(n57) );
  INV2_8TH40 U43 ( .I(B[9]), .ZN(n61) );
  INV2_8TH40 U44 ( .I(B[12]), .ZN(n34) );
  INV2_8TH40 U45 ( .I(B[16]), .ZN(n38) );
  INV2_8TH40 U46 ( .I(B[23]), .ZN(n46) );
  INV2_8TH40 U47 ( .I(B[27]), .ZN(n50) );
  INV2_8TH40 U48 ( .I(B[30]), .ZN(n54) );
  INV2_8TH40 U49 ( .I(B[3]), .ZN(n55) );
  INV2_8TH40 U50 ( .I(B[7]), .ZN(n59) );
  INV2_8TH40 U51 ( .I(B[10]), .ZN(n32) );
  INV2_8TH40 U52 ( .I(B[14]), .ZN(n36) );
  INV2_8TH40 U53 ( .I(B[18]), .ZN(n40) );
  INV2_8TH40 U54 ( .I(B[21]), .ZN(n44) );
  INV2_8TH40 U55 ( .I(B[25]), .ZN(n48) );
  INV2_8TH40 U56 ( .I(B[29]), .ZN(n52) );
  INV2_8TH40 U57 ( .I(B[6]), .ZN(n58) );
  INV2_8TH40 U58 ( .I(B[13]), .ZN(n35) );
  INV2_8TH40 U59 ( .I(B[17]), .ZN(n39) );
  INV2_8TH40 U60 ( .I(B[20]), .ZN(n43) );
  INV2_8TH40 U61 ( .I(B[24]), .ZN(n47) );
  INV2_8TH40 U62 ( .I(B[28]), .ZN(n51) );
  XOR2V2_8TH40 U63 ( .A1(n23), .A2(n54), .Z(DIFF[30]) );
  XOR2V2_8TH40 U64 ( .A1(n29), .A2(n52), .Z(DIFF[29]) );
  XOR2V2_8TH40 U65 ( .A1(n15), .A2(n51), .Z(DIFF[28]) );
  XOR2V2_8TH40 U66 ( .A1(n14), .A2(n50), .Z(DIFF[27]) );
  XOR2V2_8TH40 U67 ( .A1(n22), .A2(n49), .Z(DIFF[26]) );
  XOR2V2_8TH40 U68 ( .A1(n28), .A2(n48), .Z(DIFF[25]) );
  XOR2V2_8TH40 U69 ( .A1(n13), .A2(n47), .Z(DIFF[24]) );
  XOR2V2_8TH40 U70 ( .A1(n12), .A2(n46), .Z(DIFF[23]) );
  XOR2V2_8TH40 U71 ( .A1(n21), .A2(n45), .Z(DIFF[22]) );
  XOR2V2_8TH40 U72 ( .A1(n27), .A2(n44), .Z(DIFF[21]) );
  XOR2V2_8TH40 U73 ( .A1(n11), .A2(n43), .Z(DIFF[20]) );
  XOR2V2_8TH40 U74 ( .A1(n20), .A2(n41), .Z(DIFF[19]) );
  XOR2V2_8TH40 U75 ( .A1(n26), .A2(n40), .Z(DIFF[18]) );
  XOR2V2_8TH40 U76 ( .A1(n10), .A2(n39), .Z(DIFF[17]) );
  XOR2V2_8TH40 U77 ( .A1(n9), .A2(n38), .Z(DIFF[16]) );
  XOR2V2_8TH40 U78 ( .A1(n19), .A2(n37), .Z(DIFF[15]) );
  XOR2V2_8TH40 U79 ( .A1(n25), .A2(n36), .Z(DIFF[14]) );
  XOR2V2_8TH40 U80 ( .A1(n8), .A2(n35), .Z(DIFF[13]) );
  XOR2V2_8TH40 U81 ( .A1(n7), .A2(n34), .Z(DIFF[12]) );
  XOR2V2_8TH40 U82 ( .A1(n18), .A2(n33), .Z(DIFF[11]) );
  XOR2V2_8TH40 U83 ( .A1(n6), .A2(n32), .Z(DIFF[10]) );
  XOR2V2_8TH40 U84 ( .A1(n5), .A2(n61), .Z(DIFF[9]) );
  XOR2V2_8TH40 U85 ( .A1(n17), .A2(n60), .Z(DIFF[8]) );
  XOR2V2_8TH40 U86 ( .A1(n24), .A2(n59), .Z(DIFF[7]) );
  XOR2V2_8TH40 U87 ( .A1(n4), .A2(n58), .Z(DIFF[6]) );
  XOR2V2_8TH40 U88 ( .A1(n3), .A2(n57), .Z(DIFF[5]) );
  XOR2V2_8TH40 U89 ( .A1(n16), .A2(n56), .Z(DIFF[4]) );
  XOR2V2_8TH40 U90 ( .A1(n2), .A2(n55), .Z(DIFF[3]) );
  XOR2V2_8TH40 U91 ( .A1(n1), .A2(n53), .Z(DIFF[2]) );
  XOR2V2_8TH40 U92 ( .A1(n31), .A2(n42), .Z(DIFF[1]) );
endmodule


module div_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADH1V2C_8TH40 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADH1V2C_8TH40 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADH1V2C_8TH40 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADH1V2C_8TH40 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADH1V2C_8TH40 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADH1V2C_8TH40 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADH1V2C_8TH40 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADH1V2C_8TH40 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADH1V2C_8TH40 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADH1V2C_8TH40 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADH1V2C_8TH40 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADH1V2C_8TH40 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADH1V2C_8TH40 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADH1V2C_8TH40 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADH1V2C_8TH40 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADH1V2C_8TH40 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADH1V2C_8TH40 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADH1V2C_8TH40 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADH1V2C_8TH40 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADH1V2C_8TH40 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADH1V2C_8TH40 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADH1V2C_8TH40 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADH1V2C_8TH40 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADH1V2C_8TH40 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADH1V2C_8TH40 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADH1V2C_8TH40 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADH1V2C_8TH40 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADH1V2C_8TH40 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADH1V2C_8TH40 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADH1V2C_8TH40 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV2_8TH40 U1 ( .I(A[0]), .ZN(SUM[0]) );
  CLKXOR2V2_8TH40 U2 ( .A1(carry[31]), .A2(A[31]), .Z(SUM[31]) );
endmodule


module div_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADH1V2C_8TH40 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADH1V2C_8TH40 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADH1V2C_8TH40 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADH1V2C_8TH40 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADH1V2C_8TH40 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADH1V2C_8TH40 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADH1V2C_8TH40 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADH1V2C_8TH40 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADH1V2C_8TH40 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADH1V2C_8TH40 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADH1V2C_8TH40 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADH1V2C_8TH40 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADH1V2C_8TH40 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADH1V2C_8TH40 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADH1V2C_8TH40 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADH1V2C_8TH40 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADH1V2C_8TH40 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADH1V2C_8TH40 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADH1V2C_8TH40 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADH1V2C_8TH40 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADH1V2C_8TH40 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADH1V2C_8TH40 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADH1V2C_8TH40 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADH1V2C_8TH40 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADH1V2C_8TH40 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADH1V2C_8TH40 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADH1V2C_8TH40 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADH1V2C_8TH40 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADH1V2C_8TH40 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADH1V2C_8TH40 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2V2_8TH40 U1 ( .A1(carry[31]), .A2(A[31]), .Z(SUM[31]) );
endmodule


module div_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] DIFF;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34;
  wire   [32:1] carry;

  AD1V2C_8TH40 U2_31 ( .A(A[31]), .B(n3), .CI(carry[31]), .CO(carry[32]), .S(
        DIFF[31]) );
  AD1V2C_8TH40 U2_30 ( .A(A[30]), .B(n4), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  AD1V2C_8TH40 U2_29 ( .A(A[29]), .B(n5), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  AD1V2C_8TH40 U2_28 ( .A(A[28]), .B(n6), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  AD1V2C_8TH40 U2_27 ( .A(A[27]), .B(n7), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  AD1V2C_8TH40 U2_26 ( .A(A[26]), .B(n8), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  AD1V2C_8TH40 U2_25 ( .A(A[25]), .B(n9), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  AD1V2C_8TH40 U2_24 ( .A(A[24]), .B(n10), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  AD1V2C_8TH40 U2_23 ( .A(A[23]), .B(n11), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  AD1V2C_8TH40 U2_22 ( .A(A[22]), .B(n12), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  AD1V2C_8TH40 U2_21 ( .A(A[21]), .B(n13), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  AD1V2C_8TH40 U2_20 ( .A(A[20]), .B(n14), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  AD1V2C_8TH40 U2_19 ( .A(A[19]), .B(n15), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  AD1V2C_8TH40 U2_18 ( .A(A[18]), .B(n16), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  AD1V2C_8TH40 U2_17 ( .A(A[17]), .B(n17), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  AD1V2C_8TH40 U2_16 ( .A(A[16]), .B(n18), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  AD1V2C_8TH40 U2_15 ( .A(A[15]), .B(n19), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  AD1V2C_8TH40 U2_14 ( .A(A[14]), .B(n20), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  AD1V2C_8TH40 U2_13 ( .A(A[13]), .B(n21), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  AD1V2C_8TH40 U2_12 ( .A(A[12]), .B(n22), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  AD1V2C_8TH40 U2_11 ( .A(A[11]), .B(n23), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  AD1V2C_8TH40 U2_10 ( .A(A[10]), .B(n24), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  AD1V2C_8TH40 U2_9 ( .A(A[9]), .B(n25), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  AD1V2C_8TH40 U2_8 ( .A(A[8]), .B(n26), .CI(carry[8]), .CO(carry[9]), .S(
        DIFF[8]) );
  AD1V2C_8TH40 U2_7 ( .A(A[7]), .B(n27), .CI(carry[7]), .CO(carry[8]), .S(
        DIFF[7]) );
  AD1V2C_8TH40 U2_6 ( .A(A[6]), .B(n28), .CI(carry[6]), .CO(carry[7]), .S(
        DIFF[6]) );
  AD1V2C_8TH40 U2_5 ( .A(A[5]), .B(n29), .CI(carry[5]), .CO(carry[6]), .S(
        DIFF[5]) );
  AD1V2C_8TH40 U2_4 ( .A(A[4]), .B(n30), .CI(carry[4]), .CO(carry[5]), .S(
        DIFF[4]) );
  AD1V2C_8TH40 U2_3 ( .A(A[3]), .B(n31), .CI(carry[3]), .CO(carry[4]), .S(
        DIFF[3]) );
  AD1V2C_8TH40 U2_2 ( .A(A[2]), .B(n32), .CI(carry[2]), .CO(carry[3]), .S(
        DIFF[2]) );
  AD1V2C_8TH40 U2_1 ( .A(A[1]), .B(n33), .CI(carry[1]), .CO(carry[2]), .S(
        DIFF[1]) );
  INV2_8TH40 U1 ( .I(A[0]), .ZN(n1) );
  INV2_8TH40 U2 ( .I(carry[32]), .ZN(DIFF[32]) );
  INV2_8TH40 U3 ( .I(B[12]), .ZN(n22) );
  INV2_8TH40 U4 ( .I(B[13]), .ZN(n21) );
  INV2_8TH40 U5 ( .I(B[14]), .ZN(n20) );
  INV2_8TH40 U6 ( .I(B[15]), .ZN(n19) );
  INV2_8TH40 U7 ( .I(B[16]), .ZN(n18) );
  INV2_8TH40 U8 ( .I(B[17]), .ZN(n17) );
  INV2_8TH40 U9 ( .I(B[18]), .ZN(n16) );
  INV2_8TH40 U10 ( .I(B[19]), .ZN(n15) );
  INV2_8TH40 U11 ( .I(B[20]), .ZN(n14) );
  INV2_8TH40 U12 ( .I(B[21]), .ZN(n13) );
  INV2_8TH40 U13 ( .I(B[22]), .ZN(n12) );
  INV2_8TH40 U14 ( .I(B[23]), .ZN(n11) );
  INV2_8TH40 U15 ( .I(B[24]), .ZN(n10) );
  INV2_8TH40 U16 ( .I(B[25]), .ZN(n9) );
  INV2_8TH40 U17 ( .I(B[26]), .ZN(n8) );
  INV2_8TH40 U18 ( .I(B[27]), .ZN(n7) );
  INV2_8TH40 U19 ( .I(B[28]), .ZN(n6) );
  INV2_8TH40 U20 ( .I(B[29]), .ZN(n5) );
  INV2_8TH40 U21 ( .I(B[30]), .ZN(n4) );
  INV2_8TH40 U22 ( .I(B[2]), .ZN(n32) );
  INV2_8TH40 U23 ( .I(B[3]), .ZN(n31) );
  INV2_8TH40 U24 ( .I(B[4]), .ZN(n30) );
  INV2_8TH40 U25 ( .I(B[5]), .ZN(n29) );
  INV2_8TH40 U26 ( .I(B[6]), .ZN(n28) );
  INV2_8TH40 U27 ( .I(B[7]), .ZN(n27) );
  INV2_8TH40 U28 ( .I(B[8]), .ZN(n26) );
  INV2_8TH40 U29 ( .I(B[9]), .ZN(n25) );
  INV2_8TH40 U30 ( .I(B[10]), .ZN(n24) );
  INV2_8TH40 U31 ( .I(B[11]), .ZN(n23) );
  INV2_8TH40 U32 ( .I(B[1]), .ZN(n33) );
  NAND2V2_8TH40 U33 ( .A1(n1), .A2(B[0]), .ZN(carry[1]) );
  INV2_8TH40 U34 ( .I(B[31]), .ZN(n3) );
  INV2_8TH40 U35 ( .I(B[0]), .ZN(n34) );
  XNOR2V2_8TH40 U36 ( .A1(A[0]), .A2(n34), .ZN(DIFF[0]) );
endmodule


module div ( clk, rst, signed_div, div_opdata1, div_opdata2, div_start, 
        div_res, div_done, div_cancel_BAR );
  input [31:0] div_opdata1;
  input [31:0] div_opdata2;
  output [63:0] div_res;
  input clk, rst, signed_div, div_start, div_cancel_BAR;
  output div_done;
  wire   N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N207, N208, N209, N210, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274,
         N275, N276, N277, N278, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n4, n5, n6, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, SYNOPSYS_UNCONNECTED_1;
  wire   [64:31] dividend;
  wire   [31:0] divisor;
  wire   [32:0] div_temp;
  wire   [1:0] state;
  wire   [5:0] cnt;
  wire   [5:2] add_102_carry;

  DQV4_8TH40 state_reg_0_ ( .D(n403), .CK(clk), .Q(state[0]) );
  DQV4_8TH40 state_reg_1_ ( .D(n401), .CK(clk), .Q(state[1]) );
  DQV4_8TH40 divisor_reg_31_ ( .D(n364), .CK(clk), .Q(divisor[31]) );
  DQV4_8TH40 divisor_reg_30_ ( .D(n365), .CK(clk), .Q(divisor[30]) );
  DQV4_8TH40 divisor_reg_29_ ( .D(n366), .CK(clk), .Q(divisor[29]) );
  DQV4_8TH40 divisor_reg_28_ ( .D(n367), .CK(clk), .Q(divisor[28]) );
  DQV4_8TH40 divisor_reg_27_ ( .D(n368), .CK(clk), .Q(divisor[27]) );
  DQV4_8TH40 divisor_reg_26_ ( .D(n369), .CK(clk), .Q(divisor[26]) );
  DQV4_8TH40 divisor_reg_25_ ( .D(n370), .CK(clk), .Q(divisor[25]) );
  DQV4_8TH40 divisor_reg_24_ ( .D(n371), .CK(clk), .Q(divisor[24]) );
  DQV4_8TH40 divisor_reg_23_ ( .D(n372), .CK(clk), .Q(divisor[23]) );
  DQV4_8TH40 divisor_reg_22_ ( .D(n373), .CK(clk), .Q(divisor[22]) );
  DQV4_8TH40 divisor_reg_21_ ( .D(n374), .CK(clk), .Q(divisor[21]) );
  DQV4_8TH40 divisor_reg_20_ ( .D(n375), .CK(clk), .Q(divisor[20]) );
  DQV4_8TH40 divisor_reg_19_ ( .D(n376), .CK(clk), .Q(divisor[19]) );
  DQV4_8TH40 divisor_reg_18_ ( .D(n377), .CK(clk), .Q(divisor[18]) );
  DQV4_8TH40 divisor_reg_17_ ( .D(n378), .CK(clk), .Q(divisor[17]) );
  DQV4_8TH40 divisor_reg_16_ ( .D(n379), .CK(clk), .Q(divisor[16]) );
  DQV4_8TH40 divisor_reg_15_ ( .D(n380), .CK(clk), .Q(divisor[15]) );
  DQV4_8TH40 divisor_reg_14_ ( .D(n381), .CK(clk), .Q(divisor[14]) );
  DQV4_8TH40 divisor_reg_13_ ( .D(n382), .CK(clk), .Q(divisor[13]) );
  DQV4_8TH40 divisor_reg_12_ ( .D(n383), .CK(clk), .Q(divisor[12]) );
  DQV4_8TH40 divisor_reg_11_ ( .D(n384), .CK(clk), .Q(divisor[11]) );
  DQV4_8TH40 divisor_reg_10_ ( .D(n385), .CK(clk), .Q(divisor[10]) );
  DQV4_8TH40 divisor_reg_9_ ( .D(n386), .CK(clk), .Q(divisor[9]) );
  DQV4_8TH40 divisor_reg_8_ ( .D(n387), .CK(clk), .Q(divisor[8]) );
  DQV4_8TH40 divisor_reg_7_ ( .D(n388), .CK(clk), .Q(divisor[7]) );
  DQV4_8TH40 divisor_reg_6_ ( .D(n389), .CK(clk), .Q(divisor[6]) );
  DQV4_8TH40 divisor_reg_5_ ( .D(n390), .CK(clk), .Q(divisor[5]) );
  DQV4_8TH40 divisor_reg_4_ ( .D(n391), .CK(clk), .Q(divisor[4]) );
  DQV4_8TH40 divisor_reg_3_ ( .D(n392), .CK(clk), .Q(divisor[3]) );
  DQV4_8TH40 divisor_reg_2_ ( .D(n393), .CK(clk), .Q(divisor[2]) );
  DQV4_8TH40 divisor_reg_1_ ( .D(n394), .CK(clk), .Q(divisor[1]) );
  DQV4_8TH40 divisor_reg_0_ ( .D(n395), .CK(clk), .Q(divisor[0]) );
  DQV4_8TH40 div_done_reg ( .D(n363), .CK(clk), .Q(div_done) );
  DQV4_8TH40 cnt_reg_5_ ( .D(n402), .CK(clk), .Q(cnt[5]) );
  DQV4_8TH40 cnt_reg_0_ ( .D(n400), .CK(clk), .Q(cnt[0]) );
  DQV4_8TH40 cnt_reg_1_ ( .D(n399), .CK(clk), .Q(cnt[1]) );
  DQV4_8TH40 cnt_reg_2_ ( .D(n398), .CK(clk), .Q(cnt[2]) );
  DQV4_8TH40 cnt_reg_3_ ( .D(n397), .CK(clk), .Q(cnt[3]) );
  DQV4_8TH40 cnt_reg_4_ ( .D(n396), .CK(clk), .Q(cnt[4]) );
  DQNV4_8TH40 dividend_reg_0_ ( .D(n362), .CK(clk), .QN(n110) );
  DQV4_8TH40 div_res_reg_0_ ( .D(n297), .CK(clk), .Q(div_res[0]) );
  DQNV4_8TH40 dividend_reg_1_ ( .D(n359), .CK(clk), .QN(n109) );
  DQV4_8TH40 div_res_reg_1_ ( .D(n296), .CK(clk), .Q(div_res[1]) );
  DQNV4_8TH40 dividend_reg_2_ ( .D(n358), .CK(clk), .QN(n108) );
  DQV4_8TH40 div_res_reg_2_ ( .D(n295), .CK(clk), .Q(div_res[2]) );
  DQNV4_8TH40 dividend_reg_3_ ( .D(n357), .CK(clk), .QN(n107) );
  DQV4_8TH40 div_res_reg_3_ ( .D(n294), .CK(clk), .Q(div_res[3]) );
  DQNV4_8TH40 dividend_reg_4_ ( .D(n356), .CK(clk), .QN(n106) );
  DQV4_8TH40 div_res_reg_4_ ( .D(n293), .CK(clk), .Q(div_res[4]) );
  DQNV4_8TH40 dividend_reg_5_ ( .D(n355), .CK(clk), .QN(n105) );
  DQV4_8TH40 div_res_reg_5_ ( .D(n292), .CK(clk), .Q(div_res[5]) );
  DQNV4_8TH40 dividend_reg_6_ ( .D(n354), .CK(clk), .QN(n104) );
  DQV4_8TH40 div_res_reg_6_ ( .D(n291), .CK(clk), .Q(div_res[6]) );
  DQNV4_8TH40 dividend_reg_7_ ( .D(n353), .CK(clk), .QN(n103) );
  DQV4_8TH40 div_res_reg_7_ ( .D(n290), .CK(clk), .Q(div_res[7]) );
  DQNV4_8TH40 dividend_reg_8_ ( .D(n352), .CK(clk), .QN(n102) );
  DQV4_8TH40 div_res_reg_8_ ( .D(n289), .CK(clk), .Q(div_res[8]) );
  DQNV4_8TH40 dividend_reg_9_ ( .D(n351), .CK(clk), .QN(n101) );
  DQV4_8TH40 div_res_reg_9_ ( .D(n288), .CK(clk), .Q(div_res[9]) );
  DQNV4_8TH40 dividend_reg_10_ ( .D(n350), .CK(clk), .QN(n100) );
  DQV4_8TH40 div_res_reg_10_ ( .D(n287), .CK(clk), .Q(div_res[10]) );
  DQNV4_8TH40 dividend_reg_11_ ( .D(n349), .CK(clk), .QN(n99) );
  DQV4_8TH40 div_res_reg_11_ ( .D(n286), .CK(clk), .Q(div_res[11]) );
  DQNV4_8TH40 dividend_reg_12_ ( .D(n348), .CK(clk), .QN(n98) );
  DQV4_8TH40 div_res_reg_12_ ( .D(n285), .CK(clk), .Q(div_res[12]) );
  DQNV4_8TH40 dividend_reg_13_ ( .D(n347), .CK(clk), .QN(n97) );
  DQV4_8TH40 div_res_reg_13_ ( .D(n284), .CK(clk), .Q(div_res[13]) );
  DQNV4_8TH40 dividend_reg_14_ ( .D(n346), .CK(clk), .QN(n96) );
  DQV4_8TH40 div_res_reg_14_ ( .D(n283), .CK(clk), .Q(div_res[14]) );
  DQNV4_8TH40 dividend_reg_15_ ( .D(n345), .CK(clk), .QN(n95) );
  DQV4_8TH40 div_res_reg_15_ ( .D(n282), .CK(clk), .Q(div_res[15]) );
  DQNV4_8TH40 dividend_reg_16_ ( .D(n344), .CK(clk), .QN(n94) );
  DQV4_8TH40 div_res_reg_16_ ( .D(n281), .CK(clk), .Q(div_res[16]) );
  DQNV4_8TH40 dividend_reg_17_ ( .D(n343), .CK(clk), .QN(n93) );
  DQV4_8TH40 div_res_reg_17_ ( .D(n280), .CK(clk), .Q(div_res[17]) );
  DQNV4_8TH40 dividend_reg_18_ ( .D(n342), .CK(clk), .QN(n92) );
  DQV4_8TH40 div_res_reg_18_ ( .D(n279), .CK(clk), .Q(div_res[18]) );
  DQNV4_8TH40 dividend_reg_19_ ( .D(n341), .CK(clk), .QN(n91) );
  DQV4_8TH40 div_res_reg_19_ ( .D(n278), .CK(clk), .Q(div_res[19]) );
  DQNV4_8TH40 dividend_reg_20_ ( .D(n340), .CK(clk), .QN(n90) );
  DQV4_8TH40 div_res_reg_20_ ( .D(n277), .CK(clk), .Q(div_res[20]) );
  DQNV4_8TH40 dividend_reg_21_ ( .D(n339), .CK(clk), .QN(n89) );
  DQV4_8TH40 div_res_reg_21_ ( .D(n276), .CK(clk), .Q(div_res[21]) );
  DQNV4_8TH40 dividend_reg_22_ ( .D(n338), .CK(clk), .QN(n88) );
  DQV4_8TH40 div_res_reg_22_ ( .D(n275), .CK(clk), .Q(div_res[22]) );
  DQNV4_8TH40 dividend_reg_23_ ( .D(n337), .CK(clk), .QN(n87) );
  DQV4_8TH40 div_res_reg_23_ ( .D(n274), .CK(clk), .Q(div_res[23]) );
  DQNV4_8TH40 dividend_reg_24_ ( .D(n336), .CK(clk), .QN(n86) );
  DQV4_8TH40 div_res_reg_24_ ( .D(n273), .CK(clk), .Q(div_res[24]) );
  DQNV4_8TH40 dividend_reg_25_ ( .D(n335), .CK(clk), .QN(n85) );
  DQV4_8TH40 div_res_reg_25_ ( .D(n272), .CK(clk), .Q(div_res[25]) );
  DQNV4_8TH40 dividend_reg_26_ ( .D(n334), .CK(clk), .QN(n84) );
  DQV4_8TH40 div_res_reg_26_ ( .D(n271), .CK(clk), .Q(div_res[26]) );
  DQNV4_8TH40 dividend_reg_27_ ( .D(n333), .CK(clk), .QN(n83) );
  DQV4_8TH40 div_res_reg_27_ ( .D(n270), .CK(clk), .Q(div_res[27]) );
  DQNV4_8TH40 dividend_reg_28_ ( .D(n332), .CK(clk), .QN(n82) );
  DQV4_8TH40 div_res_reg_28_ ( .D(n269), .CK(clk), .Q(div_res[28]) );
  DQNV4_8TH40 dividend_reg_29_ ( .D(n331), .CK(clk), .QN(n81) );
  DQV4_8TH40 div_res_reg_29_ ( .D(n268), .CK(clk), .Q(div_res[29]) );
  DQNV4_8TH40 dividend_reg_30_ ( .D(n330), .CK(clk), .QN(n80) );
  DQV4_8TH40 div_res_reg_30_ ( .D(n267), .CK(clk), .Q(div_res[30]) );
  DQV4_8TH40 dividend_reg_31_ ( .D(n360), .CK(clk), .Q(dividend[31]) );
  DQV4_8TH40 div_res_reg_31_ ( .D(n266), .CK(clk), .Q(div_res[31]) );
  DQNV4_8TH40 dividend_reg_32_ ( .D(n329), .CK(clk), .QN(n38) );
  DQNV4_8TH40 dividend_reg_33_ ( .D(n328), .CK(clk), .QN(n37) );
  DQV4_8TH40 div_res_reg_32_ ( .D(n265), .CK(clk), .Q(div_res[32]) );
  DQNV4_8TH40 dividend_reg_34_ ( .D(n327), .CK(clk), .QN(n36) );
  DQV4_8TH40 div_res_reg_33_ ( .D(n264), .CK(clk), .Q(div_res[33]) );
  DQNV4_8TH40 dividend_reg_35_ ( .D(n326), .CK(clk), .QN(n35) );
  DQV4_8TH40 div_res_reg_34_ ( .D(n263), .CK(clk), .Q(div_res[34]) );
  DQNV4_8TH40 dividend_reg_36_ ( .D(n325), .CK(clk), .QN(n34) );
  DQV4_8TH40 div_res_reg_35_ ( .D(n262), .CK(clk), .Q(div_res[35]) );
  DQNV4_8TH40 dividend_reg_37_ ( .D(n324), .CK(clk), .QN(n33) );
  DQV4_8TH40 div_res_reg_36_ ( .D(n261), .CK(clk), .Q(div_res[36]) );
  DQNV4_8TH40 dividend_reg_38_ ( .D(n323), .CK(clk), .QN(n32) );
  DQV4_8TH40 div_res_reg_37_ ( .D(n260), .CK(clk), .Q(div_res[37]) );
  DQNV4_8TH40 dividend_reg_39_ ( .D(n322), .CK(clk), .QN(n31) );
  DQV4_8TH40 div_res_reg_38_ ( .D(n259), .CK(clk), .Q(div_res[38]) );
  DQNV4_8TH40 dividend_reg_40_ ( .D(n321), .CK(clk), .QN(n30) );
  DQV4_8TH40 div_res_reg_39_ ( .D(n258), .CK(clk), .Q(div_res[39]) );
  DQNV4_8TH40 dividend_reg_41_ ( .D(n320), .CK(clk), .QN(n29) );
  DQV4_8TH40 div_res_reg_40_ ( .D(n257), .CK(clk), .Q(div_res[40]) );
  DQNV4_8TH40 dividend_reg_42_ ( .D(n319), .CK(clk), .QN(n28) );
  DQV4_8TH40 div_res_reg_41_ ( .D(n256), .CK(clk), .Q(div_res[41]) );
  DQNV4_8TH40 dividend_reg_43_ ( .D(n318), .CK(clk), .QN(n27) );
  DQV4_8TH40 div_res_reg_42_ ( .D(n255), .CK(clk), .Q(div_res[42]) );
  DQNV4_8TH40 dividend_reg_44_ ( .D(n317), .CK(clk), .QN(n26) );
  DQV4_8TH40 div_res_reg_43_ ( .D(n254), .CK(clk), .Q(div_res[43]) );
  DQNV4_8TH40 dividend_reg_45_ ( .D(n316), .CK(clk), .QN(n25) );
  DQV4_8TH40 div_res_reg_44_ ( .D(n253), .CK(clk), .Q(div_res[44]) );
  DQNV4_8TH40 dividend_reg_46_ ( .D(n315), .CK(clk), .QN(n24) );
  DQV4_8TH40 div_res_reg_45_ ( .D(n252), .CK(clk), .Q(div_res[45]) );
  DQNV4_8TH40 dividend_reg_47_ ( .D(n314), .CK(clk), .QN(n23) );
  DQV4_8TH40 div_res_reg_46_ ( .D(n251), .CK(clk), .Q(div_res[46]) );
  DQNV4_8TH40 dividend_reg_48_ ( .D(n313), .CK(clk), .QN(n22) );
  DQV4_8TH40 div_res_reg_47_ ( .D(n250), .CK(clk), .Q(div_res[47]) );
  DQNV4_8TH40 dividend_reg_49_ ( .D(n312), .CK(clk), .QN(n21) );
  DQV4_8TH40 div_res_reg_48_ ( .D(n249), .CK(clk), .Q(div_res[48]) );
  DQNV4_8TH40 dividend_reg_50_ ( .D(n311), .CK(clk), .QN(n20) );
  DQV4_8TH40 div_res_reg_49_ ( .D(n248), .CK(clk), .Q(div_res[49]) );
  DQNV4_8TH40 dividend_reg_51_ ( .D(n310), .CK(clk), .QN(n19) );
  DQV4_8TH40 div_res_reg_50_ ( .D(n247), .CK(clk), .Q(div_res[50]) );
  DQNV4_8TH40 dividend_reg_52_ ( .D(n309), .CK(clk), .QN(n18) );
  DQV4_8TH40 div_res_reg_51_ ( .D(n246), .CK(clk), .Q(div_res[51]) );
  DQNV4_8TH40 dividend_reg_53_ ( .D(n308), .CK(clk), .QN(n17) );
  DQV4_8TH40 div_res_reg_52_ ( .D(n245), .CK(clk), .Q(div_res[52]) );
  DQNV4_8TH40 dividend_reg_54_ ( .D(n307), .CK(clk), .QN(n16) );
  DQV4_8TH40 div_res_reg_53_ ( .D(n244), .CK(clk), .Q(div_res[53]) );
  DQNV4_8TH40 dividend_reg_55_ ( .D(n306), .CK(clk), .QN(n15) );
  DQV4_8TH40 div_res_reg_54_ ( .D(n243), .CK(clk), .Q(div_res[54]) );
  DQNV4_8TH40 dividend_reg_56_ ( .D(n305), .CK(clk), .QN(n14) );
  DQV4_8TH40 div_res_reg_55_ ( .D(n242), .CK(clk), .Q(div_res[55]) );
  DQNV4_8TH40 dividend_reg_57_ ( .D(n304), .CK(clk), .QN(n13) );
  DQV4_8TH40 div_res_reg_56_ ( .D(n241), .CK(clk), .Q(div_res[56]) );
  DQNV4_8TH40 dividend_reg_58_ ( .D(n303), .CK(clk), .QN(n12) );
  DQV4_8TH40 div_res_reg_57_ ( .D(n240), .CK(clk), .Q(div_res[57]) );
  DQNV4_8TH40 dividend_reg_59_ ( .D(n302), .CK(clk), .QN(n11) );
  DQV4_8TH40 div_res_reg_58_ ( .D(n239), .CK(clk), .Q(div_res[58]) );
  DQNV4_8TH40 dividend_reg_60_ ( .D(n301), .CK(clk), .QN(n10) );
  DQV4_8TH40 div_res_reg_59_ ( .D(n238), .CK(clk), .Q(div_res[59]) );
  DQNV4_8TH40 dividend_reg_61_ ( .D(n300), .CK(clk), .QN(n9) );
  DQV4_8TH40 div_res_reg_60_ ( .D(n237), .CK(clk), .Q(div_res[60]) );
  DQNV4_8TH40 dividend_reg_62_ ( .D(n299), .CK(clk), .QN(n8) );
  DQV4_8TH40 div_res_reg_61_ ( .D(n236), .CK(clk), .Q(div_res[61]) );
  DQNV4_8TH40 dividend_reg_63_ ( .D(n298), .CK(clk), .QN(n7) );
  DQV4_8TH40 div_res_reg_62_ ( .D(n235), .CK(clk), .Q(div_res[62]) );
  DQV4_8TH40 dividend_reg_64_ ( .D(n361), .CK(clk), .Q(dividend[64]) );
  DQV4_8TH40 div_res_reg_63_ ( .D(n234), .CK(clk), .Q(div_res[63]) );
  div_DW01_sub_0 sub_add_59_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(div_opdata1), .CI(1'b0), .DIFF({N67, N66, N65, N64, N63, 
        N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, 
        N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36}) );
  div_DW01_sub_1 sub_add_65_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(div_opdata2), .CI(1'b0), .DIFF({N133, N132, N131, N130, 
        N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, 
        N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102}) );
  div_DW01_inc_0 add_112 ( .A({n230, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
        n30, n31, n32, n33, n34, n35, n36, n37}), .SUM({N344, N343, N342, N341, 
        N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, 
        N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, 
        N316, N315, N314, N313}) );
  div_DW01_inc_1 add_108 ( .A({n197, n80, n81, n82, n83, n84, n85, n86, n87, 
        n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
        n102, n103, n104, n105, n106, n107, n108, n109, n110}), .SUM({N278, 
        N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, 
        N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, 
        N253, N252, N251, N250, N249, N248, SYNOPSYS_UNCONNECTED_1}) );
  div_DW01_sub_2 sub_32 ( .A({1'b0, n229, n228, n227, n226, n225, n224, n223, 
        n222, n221, n220, n219, n218, n217, n216, n215, n214, n213, n212, n211, 
        n210, n209, n208, n207, n206, n205, n204, n203, n202, n201, n200, n199, 
        n198}), .B({1'b0, divisor}), .CI(1'b0), .DIFF(div_temp) );
  ADH1V2C_8TH40 add_102_U1_1_1 ( .A(cnt[1]), .B(cnt[0]), .CO(add_102_carry[2]), 
        .S(N207) );
  ADH1V2C_8TH40 add_102_U1_1_2 ( .A(cnt[2]), .B(add_102_carry[2]), .CO(
        add_102_carry[3]), .S(N208) );
  ADH1V2C_8TH40 add_102_U1_1_3 ( .A(cnt[3]), .B(add_102_carry[3]), .CO(
        add_102_carry[4]), .S(N209) );
  ADH1V2C_8TH40 add_102_U1_1_4 ( .A(cnt[4]), .B(add_102_carry[4]), .CO(
        add_102_carry[5]), .S(N210) );
  AO222V4_8TH40 U3 ( .A1(N103), .A2(n63), .B1(div_opdata2[1]), .B2(n64), .C1(
        divisor[1]), .C2(n62), .Z(n394) );
  AO222V4_8TH40 U4 ( .A1(N104), .A2(n63), .B1(div_opdata2[2]), .B2(n64), .C1(
        divisor[2]), .C2(n62), .Z(n393) );
  AO222V4_8TH40 U5 ( .A1(N105), .A2(n63), .B1(div_opdata2[3]), .B2(n64), .C1(
        divisor[3]), .C2(n62), .Z(n392) );
  AO222V4_8TH40 U6 ( .A1(N106), .A2(n63), .B1(div_opdata2[4]), .B2(n64), .C1(
        divisor[4]), .C2(n62), .Z(n391) );
  AO222V4_8TH40 U7 ( .A1(N107), .A2(n63), .B1(div_opdata2[5]), .B2(n64), .C1(
        divisor[5]), .C2(n62), .Z(n390) );
  AO222V4_8TH40 U8 ( .A1(N108), .A2(n63), .B1(div_opdata2[6]), .B2(n64), .C1(
        divisor[6]), .C2(n62), .Z(n389) );
  AO222V4_8TH40 U12 ( .A1(N109), .A2(n63), .B1(div_opdata2[7]), .B2(n64), .C1(
        divisor[7]), .C2(n62), .Z(n388) );
  AO222V4_8TH40 U13 ( .A1(N110), .A2(n63), .B1(div_opdata2[8]), .B2(n64), .C1(
        divisor[8]), .C2(n62), .Z(n387) );
  AO222V4_8TH40 U14 ( .A1(N111), .A2(n63), .B1(div_opdata2[9]), .B2(n64), .C1(
        divisor[9]), .C2(n62), .Z(n386) );
  AO222V4_8TH40 U15 ( .A1(N112), .A2(n63), .B1(div_opdata2[10]), .B2(n64), 
        .C1(divisor[10]), .C2(n62), .Z(n385) );
  AO222V4_8TH40 U16 ( .A1(N113), .A2(n63), .B1(div_opdata2[11]), .B2(n64), 
        .C1(divisor[11]), .C2(n62), .Z(n384) );
  AO222V4_8TH40 U17 ( .A1(N114), .A2(n63), .B1(div_opdata2[12]), .B2(n64), 
        .C1(divisor[12]), .C2(n62), .Z(n383) );
  AO222V4_8TH40 U18 ( .A1(N115), .A2(n63), .B1(div_opdata2[13]), .B2(n64), 
        .C1(divisor[13]), .C2(n62), .Z(n382) );
  AO222V4_8TH40 U19 ( .A1(N116), .A2(n63), .B1(div_opdata2[14]), .B2(n64), 
        .C1(divisor[14]), .C2(n62), .Z(n381) );
  AO222V4_8TH40 U20 ( .A1(N117), .A2(n63), .B1(div_opdata2[15]), .B2(n64), 
        .C1(divisor[15]), .C2(n62), .Z(n380) );
  AO222V4_8TH40 U21 ( .A1(N118), .A2(n63), .B1(div_opdata2[16]), .B2(n64), 
        .C1(divisor[16]), .C2(n62), .Z(n379) );
  AO222V4_8TH40 U22 ( .A1(N119), .A2(n63), .B1(div_opdata2[17]), .B2(n64), 
        .C1(divisor[17]), .C2(n62), .Z(n378) );
  AO222V4_8TH40 U23 ( .A1(N120), .A2(n63), .B1(div_opdata2[18]), .B2(n64), 
        .C1(divisor[18]), .C2(n62), .Z(n377) );
  AO222V4_8TH40 U24 ( .A1(N121), .A2(n63), .B1(div_opdata2[19]), .B2(n64), 
        .C1(divisor[19]), .C2(n62), .Z(n376) );
  AO222V4_8TH40 U25 ( .A1(N122), .A2(n63), .B1(div_opdata2[20]), .B2(n64), 
        .C1(divisor[20]), .C2(n62), .Z(n375) );
  AO222V4_8TH40 U26 ( .A1(N123), .A2(n63), .B1(div_opdata2[21]), .B2(n64), 
        .C1(divisor[21]), .C2(n62), .Z(n374) );
  AO222V4_8TH40 U27 ( .A1(N124), .A2(n63), .B1(div_opdata2[22]), .B2(n64), 
        .C1(divisor[22]), .C2(n62), .Z(n373) );
  AO222V4_8TH40 U28 ( .A1(N125), .A2(n63), .B1(div_opdata2[23]), .B2(n64), 
        .C1(divisor[23]), .C2(n62), .Z(n372) );
  AO222V4_8TH40 U29 ( .A1(N126), .A2(n63), .B1(div_opdata2[24]), .B2(n64), 
        .C1(divisor[24]), .C2(n62), .Z(n371) );
  AO222V4_8TH40 U30 ( .A1(N127), .A2(n63), .B1(div_opdata2[25]), .B2(n64), 
        .C1(divisor[25]), .C2(n62), .Z(n370) );
  AO222V4_8TH40 U31 ( .A1(N128), .A2(n63), .B1(div_opdata2[26]), .B2(n64), 
        .C1(divisor[26]), .C2(n62), .Z(n369) );
  AO222V4_8TH40 U32 ( .A1(N129), .A2(n63), .B1(div_opdata2[27]), .B2(n64), 
        .C1(divisor[27]), .C2(n62), .Z(n368) );
  AO222V4_8TH40 U33 ( .A1(N130), .A2(n63), .B1(div_opdata2[28]), .B2(n64), 
        .C1(divisor[28]), .C2(n62), .Z(n367) );
  AO222V4_8TH40 U34 ( .A1(N131), .A2(n63), .B1(div_opdata2[29]), .B2(n64), 
        .C1(divisor[29]), .C2(n62), .Z(n366) );
  AO222V4_8TH40 U35 ( .A1(N132), .A2(n63), .B1(div_opdata2[30]), .B2(n64), 
        .C1(divisor[30]), .C2(n62), .Z(n365) );
  AO222V4_8TH40 U36 ( .A1(N133), .A2(n63), .B1(n64), .B2(div_opdata2[31]), 
        .C1(divisor[31]), .C2(n62), .Z(n364) );
  AO22V4_8TH40 U37 ( .A1(n46), .A2(cnt[4]), .B1(N210), .B2(n47), .Z(n396) );
  AO22V4_8TH40 U38 ( .A1(n46), .A2(cnt[3]), .B1(N209), .B2(n47), .Z(n397) );
  AO22V4_8TH40 U39 ( .A1(n46), .A2(cnt[2]), .B1(N208), .B2(n47), .Z(n398) );
  AO22V4_8TH40 U40 ( .A1(n46), .A2(cnt[1]), .B1(N207), .B2(n47), .Z(n399) );
  MUX2NV2_8TH40 U41 ( .I0(n43), .I1(n44), .S(cnt[5]), .ZN(n402) );
  MUX2NV2_8TH40 U42 ( .I0(n48), .I1(n49), .S(n39), .ZN(n401) );
  AOI22V2_8TH40 U43 ( .A1(div_temp[0]), .A2(n74), .B1(N313), .B2(n75), .ZN(
        n148) );
  OAI21V2_8TH40 U44 ( .A1(n42), .A2(n143), .B(n144), .ZN(n70) );
  NAND2V2_8TH40 U45 ( .A1(n183), .A2(n184), .ZN(n40) );
  NOR4V2_8TH40 U46 ( .A1(n189), .A2(n190), .A3(n191), .A4(n192), .ZN(n183) );
  NOR4V2_8TH40 U47 ( .A1(n185), .A2(n186), .A3(n187), .A4(n188), .ZN(n184) );
  OAI21V2_8TH40 U48 ( .A1(n42), .A2(n181), .B(n144), .ZN(n72) );
  AND3V2_8TH40 U49 ( .A1(n195), .A2(n196), .A3(n51), .Z(n65) );
  NAND4V2_8TH40 U50 ( .A1(n40), .A2(n51), .A3(div_start), .A4(n182), .ZN(n62)
         );
  AOI31V2_8TH40 U51 ( .A1(n40), .A2(n51), .A3(n58), .B(n59), .ZN(n48) );
  OAI22V2_8TH40 U52 ( .A1(n147), .A2(n41), .B1(n56), .B2(n197), .ZN(n146) );
  OAI21V2_8TH40 U53 ( .A1(N67), .A2(n141), .B(div_opdata1[31]), .ZN(n147) );
  I2NOR4V2_8TH40 U54 ( .A1(cnt[5]), .A2(n194), .B1(cnt[0]), .B2(cnt[1]), .ZN(
        n179) );
  OAI221V2_8TH40 U55 ( .A1(n81), .A2(n67), .B1(n80), .B2(n70), .C(n140), .ZN(
        n330) );
  AOI222V2_8TH40 U56 ( .A1(N277), .A2(n77), .B1(N65), .B2(n78), .C1(
        div_opdata1[29]), .C2(n79), .ZN(n140) );
  OAI221V2_8TH40 U57 ( .A1(n82), .A2(n67), .B1(n81), .B2(n70), .C(n139), .ZN(
        n331) );
  AOI222V2_8TH40 U58 ( .A1(N276), .A2(n77), .B1(N64), .B2(n78), .C1(
        div_opdata1[28]), .C2(n79), .ZN(n139) );
  OAI221V2_8TH40 U59 ( .A1(n83), .A2(n67), .B1(n82), .B2(n70), .C(n138), .ZN(
        n332) );
  AOI222V2_8TH40 U60 ( .A1(N275), .A2(n77), .B1(N63), .B2(n78), .C1(
        div_opdata1[27]), .C2(n79), .ZN(n138) );
  OAI221V2_8TH40 U61 ( .A1(n84), .A2(n67), .B1(n83), .B2(n70), .C(n137), .ZN(
        n333) );
  AOI222V2_8TH40 U62 ( .A1(N274), .A2(n77), .B1(N62), .B2(n78), .C1(
        div_opdata1[26]), .C2(n79), .ZN(n137) );
  OAI221V2_8TH40 U63 ( .A1(n85), .A2(n67), .B1(n84), .B2(n70), .C(n136), .ZN(
        n334) );
  AOI222V2_8TH40 U64 ( .A1(N273), .A2(n77), .B1(N61), .B2(n78), .C1(
        div_opdata1[25]), .C2(n79), .ZN(n136) );
  OAI221V2_8TH40 U65 ( .A1(n86), .A2(n67), .B1(n85), .B2(n70), .C(n135), .ZN(
        n335) );
  AOI222V2_8TH40 U66 ( .A1(N272), .A2(n77), .B1(N60), .B2(n78), .C1(
        div_opdata1[24]), .C2(n79), .ZN(n135) );
  OAI221V2_8TH40 U67 ( .A1(n87), .A2(n67), .B1(n86), .B2(n70), .C(n134), .ZN(
        n336) );
  AOI222V2_8TH40 U68 ( .A1(N271), .A2(n77), .B1(N59), .B2(n78), .C1(
        div_opdata1[23]), .C2(n79), .ZN(n134) );
  OAI221V2_8TH40 U69 ( .A1(n88), .A2(n67), .B1(n87), .B2(n70), .C(n133), .ZN(
        n337) );
  AOI222V2_8TH40 U70 ( .A1(N270), .A2(n77), .B1(N58), .B2(n78), .C1(
        div_opdata1[22]), .C2(n79), .ZN(n133) );
  OAI221V2_8TH40 U71 ( .A1(n89), .A2(n67), .B1(n88), .B2(n70), .C(n132), .ZN(
        n338) );
  AOI222V2_8TH40 U72 ( .A1(N269), .A2(n77), .B1(N57), .B2(n78), .C1(
        div_opdata1[21]), .C2(n79), .ZN(n132) );
  OAI221V2_8TH40 U73 ( .A1(n90), .A2(n67), .B1(n89), .B2(n70), .C(n131), .ZN(
        n339) );
  AOI222V2_8TH40 U74 ( .A1(N268), .A2(n77), .B1(N56), .B2(n78), .C1(
        div_opdata1[20]), .C2(n79), .ZN(n131) );
  OAI221V2_8TH40 U75 ( .A1(n91), .A2(n67), .B1(n90), .B2(n70), .C(n130), .ZN(
        n340) );
  AOI222V2_8TH40 U76 ( .A1(N267), .A2(n77), .B1(N55), .B2(n78), .C1(
        div_opdata1[19]), .C2(n79), .ZN(n130) );
  OAI221V2_8TH40 U77 ( .A1(n92), .A2(n67), .B1(n91), .B2(n70), .C(n129), .ZN(
        n341) );
  AOI222V2_8TH40 U78 ( .A1(N266), .A2(n77), .B1(N54), .B2(n78), .C1(
        div_opdata1[18]), .C2(n79), .ZN(n129) );
  OAI221V2_8TH40 U79 ( .A1(n93), .A2(n67), .B1(n92), .B2(n70), .C(n128), .ZN(
        n342) );
  AOI222V2_8TH40 U80 ( .A1(N265), .A2(n77), .B1(N53), .B2(n78), .C1(
        div_opdata1[17]), .C2(n79), .ZN(n128) );
  OAI221V2_8TH40 U81 ( .A1(n94), .A2(n67), .B1(n93), .B2(n70), .C(n127), .ZN(
        n343) );
  AOI222V2_8TH40 U82 ( .A1(N264), .A2(n77), .B1(N52), .B2(n78), .C1(
        div_opdata1[16]), .C2(n79), .ZN(n127) );
  OAI221V2_8TH40 U83 ( .A1(n95), .A2(n67), .B1(n94), .B2(n70), .C(n126), .ZN(
        n344) );
  AOI222V2_8TH40 U84 ( .A1(N263), .A2(n77), .B1(N51), .B2(n78), .C1(
        div_opdata1[15]), .C2(n79), .ZN(n126) );
  OAI221V2_8TH40 U85 ( .A1(n96), .A2(n67), .B1(n95), .B2(n70), .C(n125), .ZN(
        n345) );
  AOI222V2_8TH40 U86 ( .A1(N262), .A2(n77), .B1(N50), .B2(n78), .C1(
        div_opdata1[14]), .C2(n79), .ZN(n125) );
  OAI221V2_8TH40 U87 ( .A1(n97), .A2(n67), .B1(n96), .B2(n70), .C(n124), .ZN(
        n346) );
  AOI222V2_8TH40 U88 ( .A1(N261), .A2(n77), .B1(N49), .B2(n78), .C1(
        div_opdata1[13]), .C2(n79), .ZN(n124) );
  OAI221V2_8TH40 U89 ( .A1(n98), .A2(n67), .B1(n97), .B2(n70), .C(n123), .ZN(
        n347) );
  AOI222V2_8TH40 U90 ( .A1(N260), .A2(n77), .B1(N48), .B2(n78), .C1(
        div_opdata1[12]), .C2(n79), .ZN(n123) );
  OAI221V2_8TH40 U91 ( .A1(n99), .A2(n67), .B1(n98), .B2(n70), .C(n122), .ZN(
        n348) );
  AOI222V2_8TH40 U92 ( .A1(N259), .A2(n77), .B1(N47), .B2(n78), .C1(
        div_opdata1[11]), .C2(n79), .ZN(n122) );
  OAI221V2_8TH40 U93 ( .A1(n100), .A2(n67), .B1(n99), .B2(n70), .C(n121), .ZN(
        n349) );
  AOI222V2_8TH40 U94 ( .A1(N258), .A2(n77), .B1(N46), .B2(n78), .C1(
        div_opdata1[10]), .C2(n79), .ZN(n121) );
  OAI221V2_8TH40 U95 ( .A1(n101), .A2(n67), .B1(n100), .B2(n70), .C(n120), 
        .ZN(n350) );
  AOI222V2_8TH40 U96 ( .A1(N257), .A2(n77), .B1(N45), .B2(n78), .C1(
        div_opdata1[9]), .C2(n79), .ZN(n120) );
  OAI221V2_8TH40 U97 ( .A1(n102), .A2(n67), .B1(n101), .B2(n70), .C(n119), 
        .ZN(n351) );
  AOI222V2_8TH40 U98 ( .A1(N256), .A2(n77), .B1(N44), .B2(n78), .C1(
        div_opdata1[8]), .C2(n79), .ZN(n119) );
  OAI221V2_8TH40 U99 ( .A1(n103), .A2(n67), .B1(n102), .B2(n70), .C(n118), 
        .ZN(n352) );
  AOI222V2_8TH40 U100 ( .A1(N255), .A2(n77), .B1(N43), .B2(n78), .C1(
        div_opdata1[7]), .C2(n79), .ZN(n118) );
  OAI221V2_8TH40 U101 ( .A1(n104), .A2(n67), .B1(n103), .B2(n70), .C(n117), 
        .ZN(n353) );
  AOI222V2_8TH40 U102 ( .A1(N254), .A2(n77), .B1(N42), .B2(n78), .C1(
        div_opdata1[6]), .C2(n79), .ZN(n117) );
  OAI221V2_8TH40 U103 ( .A1(n105), .A2(n67), .B1(n104), .B2(n70), .C(n116), 
        .ZN(n354) );
  AOI222V2_8TH40 U104 ( .A1(N253), .A2(n77), .B1(N41), .B2(n78), .C1(
        div_opdata1[5]), .C2(n79), .ZN(n116) );
  OAI221V2_8TH40 U105 ( .A1(n106), .A2(n67), .B1(n105), .B2(n70), .C(n115), 
        .ZN(n355) );
  AOI222V2_8TH40 U106 ( .A1(N252), .A2(n77), .B1(N40), .B2(n78), .C1(
        div_opdata1[4]), .C2(n79), .ZN(n115) );
  OAI221V2_8TH40 U107 ( .A1(n107), .A2(n67), .B1(n106), .B2(n70), .C(n114), 
        .ZN(n356) );
  AOI222V2_8TH40 U108 ( .A1(N251), .A2(n77), .B1(N39), .B2(n78), .C1(
        div_opdata1[3]), .C2(n79), .ZN(n114) );
  OAI221V2_8TH40 U109 ( .A1(n108), .A2(n67), .B1(n107), .B2(n70), .C(n113), 
        .ZN(n357) );
  AOI222V2_8TH40 U110 ( .A1(N250), .A2(n77), .B1(N38), .B2(n78), .C1(
        div_opdata1[2]), .C2(n79), .ZN(n113) );
  OAI221V2_8TH40 U111 ( .A1(n109), .A2(n67), .B1(n108), .B2(n70), .C(n112), 
        .ZN(n358) );
  AOI222V2_8TH40 U112 ( .A1(N249), .A2(n77), .B1(N37), .B2(n78), .C1(
        div_opdata1[1]), .C2(n79), .ZN(n112) );
  OAI221V2_8TH40 U113 ( .A1(n110), .A2(n67), .B1(n109), .B2(n70), .C(n111), 
        .ZN(n359) );
  AOI222V2_8TH40 U114 ( .A1(N248), .A2(n77), .B1(N36), .B2(n78), .C1(
        div_opdata1[0]), .C2(n79), .ZN(n111) );
  OAI221V2_8TH40 U115 ( .A1(n80), .A2(n67), .B1(n197), .B2(n70), .C(n76), .ZN(
        n360) );
  AOI222V2_8TH40 U116 ( .A1(N278), .A2(n77), .B1(N66), .B2(n78), .C1(
        div_opdata1[30]), .C2(n79), .ZN(n76) );
  OAI221V2_8TH40 U117 ( .A1(n8), .A2(n71), .B1(n7), .B2(n72), .C(n178), .ZN(
        n298) );
  AOI22V2_8TH40 U118 ( .A1(div_temp[30]), .A2(n74), .B1(N343), .B2(n75), .ZN(
        n178) );
  OAI221V2_8TH40 U119 ( .A1(n9), .A2(n71), .B1(n8), .B2(n72), .C(n177), .ZN(
        n299) );
  AOI22V2_8TH40 U120 ( .A1(div_temp[29]), .A2(n74), .B1(N342), .B2(n75), .ZN(
        n177) );
  OAI221V2_8TH40 U121 ( .A1(n10), .A2(n71), .B1(n9), .B2(n72), .C(n176), .ZN(
        n300) );
  AOI22V2_8TH40 U122 ( .A1(div_temp[28]), .A2(n74), .B1(N341), .B2(n75), .ZN(
        n176) );
  OAI221V2_8TH40 U123 ( .A1(n11), .A2(n71), .B1(n10), .B2(n72), .C(n175), .ZN(
        n301) );
  AOI22V2_8TH40 U124 ( .A1(div_temp[27]), .A2(n74), .B1(N340), .B2(n75), .ZN(
        n175) );
  OAI221V2_8TH40 U125 ( .A1(n12), .A2(n71), .B1(n11), .B2(n72), .C(n174), .ZN(
        n302) );
  AOI22V2_8TH40 U126 ( .A1(div_temp[26]), .A2(n74), .B1(N339), .B2(n75), .ZN(
        n174) );
  OAI221V2_8TH40 U127 ( .A1(n13), .A2(n71), .B1(n12), .B2(n72), .C(n173), .ZN(
        n303) );
  AOI22V2_8TH40 U128 ( .A1(div_temp[25]), .A2(n74), .B1(N338), .B2(n75), .ZN(
        n173) );
  OAI221V2_8TH40 U129 ( .A1(n14), .A2(n71), .B1(n13), .B2(n72), .C(n172), .ZN(
        n304) );
  AOI22V2_8TH40 U130 ( .A1(div_temp[24]), .A2(n74), .B1(N337), .B2(n75), .ZN(
        n172) );
  OAI221V2_8TH40 U131 ( .A1(n15), .A2(n71), .B1(n14), .B2(n72), .C(n171), .ZN(
        n305) );
  AOI22V2_8TH40 U132 ( .A1(div_temp[23]), .A2(n74), .B1(N336), .B2(n75), .ZN(
        n171) );
  OAI221V2_8TH40 U133 ( .A1(n16), .A2(n71), .B1(n15), .B2(n72), .C(n170), .ZN(
        n306) );
  AOI22V2_8TH40 U134 ( .A1(div_temp[22]), .A2(n74), .B1(N335), .B2(n75), .ZN(
        n170) );
  OAI221V2_8TH40 U135 ( .A1(n17), .A2(n71), .B1(n16), .B2(n72), .C(n169), .ZN(
        n307) );
  AOI22V2_8TH40 U136 ( .A1(div_temp[21]), .A2(n74), .B1(N334), .B2(n75), .ZN(
        n169) );
  OAI221V2_8TH40 U137 ( .A1(n18), .A2(n71), .B1(n17), .B2(n72), .C(n168), .ZN(
        n308) );
  AOI22V2_8TH40 U138 ( .A1(div_temp[20]), .A2(n74), .B1(N333), .B2(n75), .ZN(
        n168) );
  OAI221V2_8TH40 U139 ( .A1(n19), .A2(n71), .B1(n18), .B2(n72), .C(n167), .ZN(
        n309) );
  AOI22V2_8TH40 U140 ( .A1(div_temp[19]), .A2(n74), .B1(N332), .B2(n75), .ZN(
        n167) );
  OAI221V2_8TH40 U141 ( .A1(n20), .A2(n71), .B1(n19), .B2(n72), .C(n166), .ZN(
        n310) );
  AOI22V2_8TH40 U142 ( .A1(div_temp[18]), .A2(n74), .B1(N331), .B2(n75), .ZN(
        n166) );
  OAI221V2_8TH40 U143 ( .A1(n21), .A2(n71), .B1(n20), .B2(n72), .C(n165), .ZN(
        n311) );
  AOI22V2_8TH40 U144 ( .A1(div_temp[17]), .A2(n74), .B1(N330), .B2(n75), .ZN(
        n165) );
  OAI221V2_8TH40 U145 ( .A1(n22), .A2(n71), .B1(n21), .B2(n72), .C(n164), .ZN(
        n312) );
  AOI22V2_8TH40 U146 ( .A1(div_temp[16]), .A2(n74), .B1(N329), .B2(n75), .ZN(
        n164) );
  OAI221V2_8TH40 U147 ( .A1(n23), .A2(n71), .B1(n22), .B2(n72), .C(n163), .ZN(
        n313) );
  AOI22V2_8TH40 U148 ( .A1(div_temp[15]), .A2(n74), .B1(N328), .B2(n75), .ZN(
        n163) );
  OAI221V2_8TH40 U149 ( .A1(n24), .A2(n71), .B1(n23), .B2(n72), .C(n162), .ZN(
        n314) );
  AOI22V2_8TH40 U150 ( .A1(div_temp[14]), .A2(n74), .B1(N327), .B2(n75), .ZN(
        n162) );
  OAI221V2_8TH40 U151 ( .A1(n25), .A2(n71), .B1(n24), .B2(n72), .C(n161), .ZN(
        n315) );
  AOI22V2_8TH40 U152 ( .A1(div_temp[13]), .A2(n74), .B1(N326), .B2(n75), .ZN(
        n161) );
  OAI221V2_8TH40 U153 ( .A1(n26), .A2(n71), .B1(n25), .B2(n72), .C(n160), .ZN(
        n316) );
  AOI22V2_8TH40 U154 ( .A1(div_temp[12]), .A2(n74), .B1(N325), .B2(n75), .ZN(
        n160) );
  OAI221V2_8TH40 U155 ( .A1(n27), .A2(n71), .B1(n26), .B2(n72), .C(n159), .ZN(
        n317) );
  AOI22V2_8TH40 U156 ( .A1(div_temp[11]), .A2(n74), .B1(N324), .B2(n75), .ZN(
        n159) );
  OAI221V2_8TH40 U157 ( .A1(n28), .A2(n71), .B1(n27), .B2(n72), .C(n158), .ZN(
        n318) );
  AOI22V2_8TH40 U158 ( .A1(div_temp[10]), .A2(n74), .B1(N323), .B2(n75), .ZN(
        n158) );
  OAI221V2_8TH40 U159 ( .A1(n29), .A2(n71), .B1(n28), .B2(n72), .C(n157), .ZN(
        n319) );
  AOI22V2_8TH40 U160 ( .A1(div_temp[9]), .A2(n74), .B1(N322), .B2(n75), .ZN(
        n157) );
  OAI221V2_8TH40 U161 ( .A1(n30), .A2(n71), .B1(n29), .B2(n72), .C(n156), .ZN(
        n320) );
  AOI22V2_8TH40 U162 ( .A1(div_temp[8]), .A2(n74), .B1(N321), .B2(n75), .ZN(
        n156) );
  OAI221V2_8TH40 U163 ( .A1(n31), .A2(n71), .B1(n30), .B2(n72), .C(n155), .ZN(
        n321) );
  AOI22V2_8TH40 U164 ( .A1(div_temp[7]), .A2(n74), .B1(N320), .B2(n75), .ZN(
        n155) );
  OAI221V2_8TH40 U165 ( .A1(n32), .A2(n71), .B1(n31), .B2(n72), .C(n154), .ZN(
        n322) );
  AOI22V2_8TH40 U166 ( .A1(div_temp[6]), .A2(n74), .B1(N319), .B2(n75), .ZN(
        n154) );
  OAI221V2_8TH40 U167 ( .A1(n33), .A2(n71), .B1(n32), .B2(n72), .C(n153), .ZN(
        n323) );
  AOI22V2_8TH40 U168 ( .A1(div_temp[5]), .A2(n74), .B1(N318), .B2(n75), .ZN(
        n153) );
  OAI221V2_8TH40 U169 ( .A1(n34), .A2(n71), .B1(n33), .B2(n72), .C(n152), .ZN(
        n324) );
  AOI22V2_8TH40 U170 ( .A1(div_temp[4]), .A2(n74), .B1(N317), .B2(n75), .ZN(
        n152) );
  OAI221V2_8TH40 U171 ( .A1(n35), .A2(n71), .B1(n34), .B2(n72), .C(n151), .ZN(
        n325) );
  AOI22V2_8TH40 U172 ( .A1(div_temp[3]), .A2(n74), .B1(N316), .B2(n75), .ZN(
        n151) );
  OAI221V2_8TH40 U173 ( .A1(n36), .A2(n71), .B1(n35), .B2(n72), .C(n150), .ZN(
        n326) );
  AOI22V2_8TH40 U174 ( .A1(div_temp[2]), .A2(n74), .B1(N315), .B2(n75), .ZN(
        n150) );
  OAI221V2_8TH40 U175 ( .A1(n37), .A2(n71), .B1(n36), .B2(n72), .C(n149), .ZN(
        n327) );
  AOI22V2_8TH40 U176 ( .A1(div_temp[1]), .A2(n74), .B1(N314), .B2(n75), .ZN(
        n149) );
  OAI221V2_8TH40 U177 ( .A1(n7), .A2(n71), .B1(n230), .B2(n72), .C(n73), .ZN(
        n361) );
  AOI22V2_8TH40 U178 ( .A1(div_temp[31]), .A2(n74), .B1(N344), .B2(n75), .ZN(
        n73) );
  OAI21V2_8TH40 U179 ( .A1(div_temp[32]), .A2(n67), .B(n68), .ZN(n362) );
  I2NOR3V2_8TH40 U180 ( .A1(n50), .A2(n51), .B(n52), .ZN(n39) );
  OAOI211V2_8TH40 U181 ( .A1(n49), .A2(n53), .B(state[0]), .C(n54), .ZN(n50)
         );
  INV2_8TH40 U182 ( .I(dividend[64]), .ZN(n230) );
  INV2_8TH40 U183 ( .I(dividend[31]), .ZN(n197) );
  NAND2V2_8TH40 U184 ( .A1(n4), .A2(n5), .ZN(n403) );
  CLKNV1_8TH40 U185 ( .I(n37), .ZN(n199) );
  CLKNV1_8TH40 U186 ( .I(n36), .ZN(n200) );
  CLKNV1_8TH40 U187 ( .I(n35), .ZN(n201) );
  CLKNV1_8TH40 U188 ( .I(n34), .ZN(n202) );
  CLKNV1_8TH40 U189 ( .I(n33), .ZN(n203) );
  CLKNV1_8TH40 U190 ( .I(n32), .ZN(n204) );
  CLKNV1_8TH40 U191 ( .I(n31), .ZN(n205) );
  CLKNV1_8TH40 U192 ( .I(n30), .ZN(n206) );
  CLKNV1_8TH40 U193 ( .I(n29), .ZN(n207) );
  CLKNV1_8TH40 U194 ( .I(n28), .ZN(n208) );
  CLKNV1_8TH40 U195 ( .I(n27), .ZN(n209) );
  CLKNV1_8TH40 U196 ( .I(n26), .ZN(n210) );
  CLKNV1_8TH40 U197 ( .I(n25), .ZN(n211) );
  CLKNV1_8TH40 U198 ( .I(n24), .ZN(n212) );
  CLKNV1_8TH40 U199 ( .I(n23), .ZN(n213) );
  CLKNV1_8TH40 U200 ( .I(n22), .ZN(n214) );
  CLKNV1_8TH40 U201 ( .I(n21), .ZN(n215) );
  CLKNV1_8TH40 U202 ( .I(n20), .ZN(n216) );
  CLKNV1_8TH40 U203 ( .I(n19), .ZN(n217) );
  CLKNV1_8TH40 U204 ( .I(n18), .ZN(n218) );
  CLKNV1_8TH40 U205 ( .I(n17), .ZN(n219) );
  CLKNV1_8TH40 U206 ( .I(n16), .ZN(n220) );
  CLKNV1_8TH40 U207 ( .I(n15), .ZN(n221) );
  CLKNV1_8TH40 U208 ( .I(n14), .ZN(n222) );
  CLKNV1_8TH40 U209 ( .I(n13), .ZN(n223) );
  CLKNV1_8TH40 U210 ( .I(n12), .ZN(n224) );
  CLKNV1_8TH40 U211 ( .I(n11), .ZN(n225) );
  CLKNV1_8TH40 U212 ( .I(n10), .ZN(n226) );
  CLKNV1_8TH40 U213 ( .I(n9), .ZN(n227) );
  CLKNV1_8TH40 U214 ( .I(n8), .ZN(n228) );
  CLKNV1_8TH40 U215 ( .I(n7), .ZN(n229) );
  MUX2NV0_8TH40 U216 ( .I0(n6), .I1(state[0]), .S(n39), .ZN(n4) );
  OAI31V0_8TH40 U217 ( .A1(n40), .A2(rst), .A3(n41), .B(n42), .ZN(n6) );
  IAO21V0_8TH40 U218 ( .A1(n45), .A2(add_102_carry[5]), .B(n46), .ZN(n44) );
  CLKNAND2V1_8TH40 U219 ( .A1(add_102_carry[5]), .A2(n47), .ZN(n43) );
  MUX2NV0_8TH40 U220 ( .I0(n55), .I1(n56), .S(n57), .ZN(n54) );
  CLKNAND2V1_8TH40 U221 ( .A1(n58), .A2(div_start), .ZN(n55) );
  CLKNAND2V1_8TH40 U222 ( .A1(n42), .A2(n5), .ZN(n59) );
  MUX2NV0_8TH40 U223 ( .I0(n45), .I1(n60), .S(cnt[0]), .ZN(n400) );
  CLKNV1_8TH40 U224 ( .I(n45), .ZN(n47) );
  CLKNAND2V1_8TH40 U225 ( .A1(n61), .A2(n60), .ZN(n45) );
  CLKNV1_8TH40 U226 ( .I(n60), .ZN(n46) );
  CLKNAND2V1_8TH40 U227 ( .A1(n62), .A2(n42), .ZN(n60) );
  AO222V0_8TH40 U228 ( .A1(N102), .A2(n63), .B1(div_opdata2[0]), .B2(n64), 
        .C1(divisor[0]), .C2(n62), .Z(n395) );
  AOI21V0_8TH40 U229 ( .A1(div_opdata2[31]), .A2(signed_div), .B(n62), .ZN(n64) );
  I2NOR3V1_8TH40 U230 ( .A1(div_opdata2[31]), .A2(signed_div), .B(n62), .ZN(
        n63) );
  IOA21V0_8TH40 U231 ( .A1(div_done), .A2(n65), .B(n66), .ZN(n363) );
  AO21V0_8TH40 U232 ( .A1(n69), .A2(n70), .B(n110), .Z(n68) );
  AND3V0_8TH40 U233 ( .A1(n70), .A2(n141), .A3(n58), .Z(n79) );
  AND3V0_8TH40 U234 ( .A1(n58), .A2(n70), .A3(n142), .Z(n78) );
  CLKNV1_8TH40 U235 ( .I(n69), .ZN(n77) );
  CLKNAND2V1_8TH40 U236 ( .A1(n52), .A2(n70), .ZN(n69) );
  CLKNAND2V1_8TH40 U237 ( .A1(n61), .A2(n70), .ZN(n67) );
  MUX2NV0_8TH40 U238 ( .I0(n142), .I1(n145), .S(div_opdata2[31]), .ZN(n143) );
  CKMUX2V2_8TH40 U239 ( .I0(n146), .I1(n198), .S(n144), .Z(n329) );
  CLKNV1_8TH40 U240 ( .I(n38), .ZN(n198) );
  OAI221V0_8TH40 U241 ( .A1(n38), .A2(n71), .B1(n37), .B2(n72), .C(n148), .ZN(
        n328) );
  AND2V0_8TH40 U242 ( .A1(n52), .A2(n72), .Z(n75) );
  AND2V0_8TH40 U243 ( .A1(n179), .A2(n180), .Z(n52) );
  I2NOR3V1_8TH40 U244 ( .A1(n72), .A2(n61), .B(div_temp[32]), .ZN(n74) );
  NAND3V0P5_8TH40 U245 ( .A1(n61), .A2(n72), .A3(div_temp[32]), .ZN(n71) );
  OA211V0_8TH40 U246 ( .A1(n179), .A2(n42), .B(n62), .C(n5), .Z(n144) );
  NAND3V0P5_8TH40 U247 ( .A1(n51), .A2(n49), .A3(state[0]), .ZN(n5) );
  NOR2V0P5_8TH40 U248 ( .A1(n41), .A2(n57), .ZN(n182) );
  CLKNV1_8TH40 U249 ( .I(n58), .ZN(n41) );
  OR4V0_8TH40 U250 ( .A1(div_opdata2[24]), .A2(div_opdata2[25]), .A3(
        div_opdata2[26]), .A4(div_opdata2[27]), .Z(n188) );
  OR4V0_8TH40 U251 ( .A1(div_opdata2[28]), .A2(div_opdata2[29]), .A3(
        div_opdata2[2]), .A4(div_opdata2[30]), .Z(n187) );
  OR4V0_8TH40 U252 ( .A1(div_opdata2[31]), .A2(div_opdata2[3]), .A3(
        div_opdata2[4]), .A4(div_opdata2[5]), .Z(n186) );
  OR4V0_8TH40 U253 ( .A1(div_opdata2[6]), .A2(div_opdata2[7]), .A3(
        div_opdata2[8]), .A4(div_opdata2[9]), .Z(n185) );
  OR4V0_8TH40 U254 ( .A1(div_opdata2[0]), .A2(div_opdata2[10]), .A3(
        div_opdata2[11]), .A4(div_opdata2[12]), .Z(n192) );
  OR4V0_8TH40 U255 ( .A1(div_opdata2[13]), .A2(div_opdata2[14]), .A3(
        div_opdata2[15]), .A4(div_opdata2[16]), .Z(n191) );
  OR4V0_8TH40 U256 ( .A1(div_opdata2[17]), .A2(div_opdata2[18]), .A3(
        div_opdata2[19]), .A4(div_opdata2[1]), .Z(n190) );
  OR4V0_8TH40 U257 ( .A1(div_opdata2[20]), .A2(div_opdata2[21]), .A3(
        div_opdata2[22]), .A4(div_opdata2[23]), .Z(n189) );
  MUX2NV0_8TH40 U258 ( .I0(n145), .I1(n142), .S(n230), .ZN(n181) );
  CLKNV1_8TH40 U259 ( .I(n141), .ZN(n142) );
  CLKNAND2V1_8TH40 U260 ( .A1(signed_div), .A2(div_opdata1[31]), .ZN(n141) );
  NOR2V0P5_8TH40 U261 ( .A1(div_opdata1[31]), .A2(n193), .ZN(n145) );
  CLKNV1_8TH40 U262 ( .I(signed_div), .ZN(n193) );
  NAND3V0P5_8TH40 U263 ( .A1(n180), .A2(n51), .A3(div_cancel_BAR), .ZN(n42) );
  NOR2V0P5_8TH40 U264 ( .A1(n56), .A2(n179), .ZN(n61) );
  NOR3V0P5_8TH40 U265 ( .A1(cnt[2]), .A2(cnt[4]), .A3(cnt[3]), .ZN(n194) );
  CLKNV1_8TH40 U266 ( .I(n180), .ZN(n56) );
  NOR2V0P5_8TH40 U267 ( .A1(n49), .A2(state[0]), .ZN(n180) );
  CLKNV1_8TH40 U268 ( .I(state[1]), .ZN(n49) );
  IOA22V0_8TH40 U269 ( .B1(n110), .B2(n66), .A1(div_res[0]), .A2(n65), .ZN(
        n297) );
  IOA22V0_8TH40 U270 ( .B1(n109), .B2(n66), .A1(div_res[1]), .A2(n65), .ZN(
        n296) );
  IOA22V0_8TH40 U271 ( .B1(n108), .B2(n66), .A1(div_res[2]), .A2(n65), .ZN(
        n295) );
  IOA22V0_8TH40 U272 ( .B1(n107), .B2(n66), .A1(div_res[3]), .A2(n65), .ZN(
        n294) );
  IOA22V0_8TH40 U273 ( .B1(n106), .B2(n66), .A1(div_res[4]), .A2(n65), .ZN(
        n293) );
  IOA22V0_8TH40 U274 ( .B1(n105), .B2(n66), .A1(div_res[5]), .A2(n65), .ZN(
        n292) );
  IOA22V0_8TH40 U275 ( .B1(n104), .B2(n66), .A1(div_res[6]), .A2(n65), .ZN(
        n291) );
  IOA22V0_8TH40 U276 ( .B1(n103), .B2(n66), .A1(div_res[7]), .A2(n65), .ZN(
        n290) );
  IOA22V0_8TH40 U277 ( .B1(n102), .B2(n66), .A1(div_res[8]), .A2(n65), .ZN(
        n289) );
  IOA22V0_8TH40 U278 ( .B1(n101), .B2(n66), .A1(div_res[9]), .A2(n65), .ZN(
        n288) );
  IOA22V0_8TH40 U279 ( .B1(n100), .B2(n66), .A1(div_res[10]), .A2(n65), .ZN(
        n287) );
  IOA22V0_8TH40 U280 ( .B1(n99), .B2(n66), .A1(div_res[11]), .A2(n65), .ZN(
        n286) );
  IOA22V0_8TH40 U281 ( .B1(n98), .B2(n66), .A1(div_res[12]), .A2(n65), .ZN(
        n285) );
  IOA22V0_8TH40 U282 ( .B1(n97), .B2(n66), .A1(div_res[13]), .A2(n65), .ZN(
        n284) );
  IOA22V0_8TH40 U283 ( .B1(n96), .B2(n66), .A1(div_res[14]), .A2(n65), .ZN(
        n283) );
  IOA22V0_8TH40 U284 ( .B1(n95), .B2(n66), .A1(div_res[15]), .A2(n65), .ZN(
        n282) );
  IOA22V0_8TH40 U285 ( .B1(n94), .B2(n66), .A1(div_res[16]), .A2(n65), .ZN(
        n281) );
  IOA22V0_8TH40 U286 ( .B1(n93), .B2(n66), .A1(div_res[17]), .A2(n65), .ZN(
        n280) );
  IOA22V0_8TH40 U287 ( .B1(n92), .B2(n66), .A1(div_res[18]), .A2(n65), .ZN(
        n279) );
  IOA22V0_8TH40 U288 ( .B1(n91), .B2(n66), .A1(div_res[19]), .A2(n65), .ZN(
        n278) );
  IOA22V0_8TH40 U289 ( .B1(n90), .B2(n66), .A1(div_res[20]), .A2(n65), .ZN(
        n277) );
  IOA22V0_8TH40 U290 ( .B1(n89), .B2(n66), .A1(div_res[21]), .A2(n65), .ZN(
        n276) );
  IOA22V0_8TH40 U291 ( .B1(n88), .B2(n66), .A1(div_res[22]), .A2(n65), .ZN(
        n275) );
  IOA22V0_8TH40 U292 ( .B1(n87), .B2(n66), .A1(div_res[23]), .A2(n65), .ZN(
        n274) );
  IOA22V0_8TH40 U293 ( .B1(n86), .B2(n66), .A1(div_res[24]), .A2(n65), .ZN(
        n273) );
  IOA22V0_8TH40 U294 ( .B1(n85), .B2(n66), .A1(div_res[25]), .A2(n65), .ZN(
        n272) );
  IOA22V0_8TH40 U295 ( .B1(n84), .B2(n66), .A1(div_res[26]), .A2(n65), .ZN(
        n271) );
  IOA22V0_8TH40 U296 ( .B1(n83), .B2(n66), .A1(div_res[27]), .A2(n65), .ZN(
        n270) );
  IOA22V0_8TH40 U297 ( .B1(n82), .B2(n66), .A1(div_res[28]), .A2(n65), .ZN(
        n269) );
  IOA22V0_8TH40 U298 ( .B1(n81), .B2(n66), .A1(div_res[29]), .A2(n65), .ZN(
        n268) );
  IOA22V0_8TH40 U299 ( .B1(n80), .B2(n66), .A1(div_res[30]), .A2(n65), .ZN(
        n267) );
  IOA22V0_8TH40 U300 ( .B1(n197), .B2(n66), .A1(div_res[31]), .A2(n65), .ZN(
        n266) );
  IOA22V0_8TH40 U301 ( .B1(n37), .B2(n66), .A1(div_res[32]), .A2(n65), .ZN(
        n265) );
  IOA22V0_8TH40 U302 ( .B1(n36), .B2(n66), .A1(div_res[33]), .A2(n65), .ZN(
        n264) );
  IOA22V0_8TH40 U303 ( .B1(n35), .B2(n66), .A1(div_res[34]), .A2(n65), .ZN(
        n263) );
  IOA22V0_8TH40 U304 ( .B1(n34), .B2(n66), .A1(div_res[35]), .A2(n65), .ZN(
        n262) );
  IOA22V0_8TH40 U305 ( .B1(n33), .B2(n66), .A1(div_res[36]), .A2(n65), .ZN(
        n261) );
  IOA22V0_8TH40 U306 ( .B1(n32), .B2(n66), .A1(div_res[37]), .A2(n65), .ZN(
        n260) );
  IOA22V0_8TH40 U307 ( .B1(n31), .B2(n66), .A1(div_res[38]), .A2(n65), .ZN(
        n259) );
  IOA22V0_8TH40 U308 ( .B1(n30), .B2(n66), .A1(div_res[39]), .A2(n65), .ZN(
        n258) );
  IOA22V0_8TH40 U309 ( .B1(n29), .B2(n66), .A1(div_res[40]), .A2(n65), .ZN(
        n257) );
  IOA22V0_8TH40 U310 ( .B1(n28), .B2(n66), .A1(div_res[41]), .A2(n65), .ZN(
        n256) );
  IOA22V0_8TH40 U311 ( .B1(n27), .B2(n66), .A1(div_res[42]), .A2(n65), .ZN(
        n255) );
  IOA22V0_8TH40 U312 ( .B1(n26), .B2(n66), .A1(div_res[43]), .A2(n65), .ZN(
        n254) );
  IOA22V0_8TH40 U313 ( .B1(n25), .B2(n66), .A1(div_res[44]), .A2(n65), .ZN(
        n253) );
  IOA22V0_8TH40 U314 ( .B1(n24), .B2(n66), .A1(div_res[45]), .A2(n65), .ZN(
        n252) );
  IOA22V0_8TH40 U315 ( .B1(n23), .B2(n66), .A1(div_res[46]), .A2(n65), .ZN(
        n251) );
  IOA22V0_8TH40 U316 ( .B1(n22), .B2(n66), .A1(div_res[47]), .A2(n65), .ZN(
        n250) );
  IOA22V0_8TH40 U317 ( .B1(n21), .B2(n66), .A1(div_res[48]), .A2(n65), .ZN(
        n249) );
  IOA22V0_8TH40 U318 ( .B1(n20), .B2(n66), .A1(div_res[49]), .A2(n65), .ZN(
        n248) );
  IOA22V0_8TH40 U319 ( .B1(n19), .B2(n66), .A1(div_res[50]), .A2(n65), .ZN(
        n247) );
  IOA22V0_8TH40 U320 ( .B1(n18), .B2(n66), .A1(div_res[51]), .A2(n65), .ZN(
        n246) );
  IOA22V0_8TH40 U321 ( .B1(n17), .B2(n66), .A1(div_res[52]), .A2(n65), .ZN(
        n245) );
  IOA22V0_8TH40 U322 ( .B1(n16), .B2(n66), .A1(div_res[53]), .A2(n65), .ZN(
        n244) );
  IOA22V0_8TH40 U323 ( .B1(n15), .B2(n66), .A1(div_res[54]), .A2(n65), .ZN(
        n243) );
  IOA22V0_8TH40 U324 ( .B1(n14), .B2(n66), .A1(div_res[55]), .A2(n65), .ZN(
        n242) );
  IOA22V0_8TH40 U325 ( .B1(n13), .B2(n66), .A1(div_res[56]), .A2(n65), .ZN(
        n241) );
  IOA22V0_8TH40 U326 ( .B1(n12), .B2(n66), .A1(div_res[57]), .A2(n65), .ZN(
        n240) );
  IOA22V0_8TH40 U327 ( .B1(n11), .B2(n66), .A1(div_res[58]), .A2(n65), .ZN(
        n239) );
  IOA22V0_8TH40 U328 ( .B1(n10), .B2(n66), .A1(div_res[59]), .A2(n65), .ZN(
        n238) );
  IOA22V0_8TH40 U329 ( .B1(n9), .B2(n66), .A1(div_res[60]), .A2(n65), .ZN(n237) );
  IOA22V0_8TH40 U330 ( .B1(n8), .B2(n66), .A1(div_res[61]), .A2(n65), .ZN(n236) );
  IOA22V0_8TH40 U331 ( .B1(n7), .B2(n66), .A1(div_res[62]), .A2(n65), .ZN(n235) );
  IOA22V0_8TH40 U332 ( .B1(n230), .B2(n66), .A1(div_res[63]), .A2(n65), .ZN(
        n234) );
  OAI21V0_8TH40 U333 ( .A1(n53), .A2(n57), .B(n58), .ZN(n196) );
  NOR2V0P5_8TH40 U334 ( .A1(state[1]), .A2(state[0]), .ZN(n58) );
  CLKNV1_8TH40 U335 ( .I(div_cancel_BAR), .ZN(n57) );
  CLKNV1_8TH40 U336 ( .I(div_start), .ZN(n53) );
  INAND3V0_8TH40 U337 ( .A1(n195), .B1(div_start), .B2(n51), .ZN(n66) );
  CLKNV1_8TH40 U338 ( .I(rst), .ZN(n51) );
  CLKNAND2V1_8TH40 U339 ( .A1(state[1]), .A2(state[0]), .ZN(n195) );
endmodule


module coprocessor0_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NOR4V2_8TH40 U1 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(EQ) );
  NAND2V2_8TH40 U2 ( .A1(n17), .A2(n18), .ZN(n4) );
  NAND4V2_8TH40 U3 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n6) );
  NAND4V2_8TH40 U4 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .ZN(n5) );
  NAND4V2_8TH40 U5 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(n3) );
  NOR4V2_8TH40 U6 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(n28) );
  NOR4V2_8TH40 U7 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(n30) );
  NOR4V2_8TH40 U8 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(n29) );
  NOR4V2_8TH40 U9 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(n18) );
  NOR4V2_8TH40 U10 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(n17) );
  NOR4V2_8TH40 U11 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(n27) );
  INV2_8TH40 U12 ( .I(B[1]), .ZN(n2) );
  INV2_8TH40 U13 ( .I(A[1]), .ZN(n1) );
  XNOR2V0_8TH40 U14 ( .A1(B[3]), .A2(A[3]), .ZN(n10) );
  XNOR2V0_8TH40 U15 ( .A1(B[4]), .A2(A[4]), .ZN(n9) );
  XNOR2V0_8TH40 U16 ( .A1(B[5]), .A2(A[5]), .ZN(n8) );
  XNOR2V0_8TH40 U17 ( .A1(B[6]), .A2(A[6]), .ZN(n7) );
  OAI22V0_8TH40 U18 ( .A1(n15), .A2(n1), .B1(B[1]), .B2(n15), .ZN(n14) );
  INOR2V0_8TH40 U19 ( .A1(B[0]), .B1(A[0]), .ZN(n15) );
  OAI22V0_8TH40 U20 ( .A1(A[1]), .A2(n16), .B1(n16), .B2(n2), .ZN(n13) );
  INOR2V0_8TH40 U21 ( .A1(A[0]), .B1(B[0]), .ZN(n16) );
  XNOR2V0_8TH40 U22 ( .A1(B[31]), .A2(A[31]), .ZN(n12) );
  XNOR2V0_8TH40 U23 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  CLKXOR2V2_8TH40 U24 ( .A1(B[10]), .A2(A[10]), .Z(n22) );
  CLKXOR2V2_8TH40 U25 ( .A1(B[9]), .A2(A[9]), .Z(n21) );
  CLKXOR2V2_8TH40 U26 ( .A1(B[8]), .A2(A[8]), .Z(n20) );
  CLKXOR2V2_8TH40 U27 ( .A1(B[7]), .A2(A[7]), .Z(n19) );
  CLKXOR2V2_8TH40 U28 ( .A1(B[14]), .A2(A[14]), .Z(n26) );
  CLKXOR2V2_8TH40 U29 ( .A1(B[13]), .A2(A[13]), .Z(n25) );
  CLKXOR2V2_8TH40 U30 ( .A1(B[12]), .A2(A[12]), .Z(n24) );
  CLKXOR2V2_8TH40 U31 ( .A1(B[11]), .A2(A[11]), .Z(n23) );
  CLKXOR2V2_8TH40 U32 ( .A1(B[18]), .A2(A[18]), .Z(n34) );
  CLKXOR2V2_8TH40 U33 ( .A1(B[17]), .A2(A[17]), .Z(n33) );
  CLKXOR2V2_8TH40 U34 ( .A1(B[16]), .A2(A[16]), .Z(n32) );
  CLKXOR2V2_8TH40 U35 ( .A1(B[15]), .A2(A[15]), .Z(n31) );
  CLKXOR2V2_8TH40 U36 ( .A1(B[22]), .A2(A[22]), .Z(n38) );
  CLKXOR2V2_8TH40 U37 ( .A1(B[21]), .A2(A[21]), .Z(n37) );
  CLKXOR2V2_8TH40 U38 ( .A1(B[20]), .A2(A[20]), .Z(n36) );
  CLKXOR2V2_8TH40 U39 ( .A1(B[19]), .A2(A[19]), .Z(n35) );
  CLKXOR2V2_8TH40 U40 ( .A1(B[26]), .A2(A[26]), .Z(n42) );
  CLKXOR2V2_8TH40 U41 ( .A1(B[25]), .A2(A[25]), .Z(n41) );
  CLKXOR2V2_8TH40 U42 ( .A1(B[24]), .A2(A[24]), .Z(n40) );
  CLKXOR2V2_8TH40 U43 ( .A1(B[23]), .A2(A[23]), .Z(n39) );
  CLKXOR2V2_8TH40 U44 ( .A1(B[30]), .A2(A[30]), .Z(n46) );
  CLKXOR2V2_8TH40 U45 ( .A1(B[29]), .A2(A[29]), .Z(n45) );
  CLKXOR2V2_8TH40 U46 ( .A1(B[28]), .A2(A[28]), .Z(n44) );
  CLKXOR2V2_8TH40 U47 ( .A1(B[27]), .A2(A[27]), .Z(n43) );
endmodule


module coprocessor0_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADH1V2C_8TH40 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADH1V2C_8TH40 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADH1V2C_8TH40 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADH1V2C_8TH40 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADH1V2C_8TH40 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADH1V2C_8TH40 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADH1V2C_8TH40 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADH1V2C_8TH40 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADH1V2C_8TH40 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADH1V2C_8TH40 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADH1V2C_8TH40 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADH1V2C_8TH40 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADH1V2C_8TH40 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADH1V2C_8TH40 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADH1V2C_8TH40 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADH1V2C_8TH40 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADH1V2C_8TH40 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADH1V2C_8TH40 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADH1V2C_8TH40 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADH1V2C_8TH40 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADH1V2C_8TH40 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADH1V2C_8TH40 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADH1V2C_8TH40 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADH1V2C_8TH40 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADH1V2C_8TH40 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADH1V2C_8TH40 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADH1V2C_8TH40 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADH1V2C_8TH40 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADH1V2C_8TH40 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADH1V2C_8TH40 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV2_8TH40 U1 ( .I(A[0]), .ZN(SUM[0]) );
  CLKXOR2V2_8TH40 U2 ( .A1(carry[31]), .A2(A[31]), .Z(SUM[31]) );
endmodule


module coprocessor0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [31:3] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = A[0];

  INV2_8TH40 U1 ( .I(carry[30]), .ZN(n1) );
  NAND2V2_8TH40 U2 ( .A1(n1), .A2(n2), .ZN(carry[31]) );
  INV2_8TH40 U3 ( .I(A[30]), .ZN(n2) );
  OR2V2_8TH40 U4 ( .A1(carry[3]), .A2(A[3]), .Z(carry[4]) );
  OR2V2_8TH40 U5 ( .A1(carry[4]), .A2(A[4]), .Z(carry[5]) );
  OR2V2_8TH40 U6 ( .A1(carry[5]), .A2(A[5]), .Z(carry[6]) );
  OR2V2_8TH40 U7 ( .A1(carry[6]), .A2(A[6]), .Z(carry[7]) );
  OR2V2_8TH40 U8 ( .A1(carry[7]), .A2(A[7]), .Z(carry[8]) );
  OR2V2_8TH40 U9 ( .A1(carry[9]), .A2(A[9]), .Z(carry[10]) );
  OR2V2_8TH40 U10 ( .A1(carry[13]), .A2(A[13]), .Z(carry[14]) );
  OR2V2_8TH40 U11 ( .A1(carry[16]), .A2(A[16]), .Z(carry[17]) );
  OR2V2_8TH40 U12 ( .A1(carry[17]), .A2(A[17]), .Z(carry[18]) );
  OR2V2_8TH40 U13 ( .A1(carry[20]), .A2(A[20]), .Z(carry[21]) );
  OR2V2_8TH40 U14 ( .A1(carry[8]), .A2(A[8]), .Z(carry[9]) );
  OR2V2_8TH40 U15 ( .A1(carry[10]), .A2(A[10]), .Z(carry[11]) );
  OR2V2_8TH40 U16 ( .A1(carry[11]), .A2(A[11]), .Z(carry[12]) );
  OR2V2_8TH40 U17 ( .A1(carry[12]), .A2(A[12]), .Z(carry[13]) );
  OR2V2_8TH40 U18 ( .A1(carry[14]), .A2(A[14]), .Z(carry[15]) );
  OR2V2_8TH40 U19 ( .A1(carry[18]), .A2(A[18]), .Z(carry[19]) );
  OR2V2_8TH40 U20 ( .A1(carry[19]), .A2(A[19]), .Z(carry[20]) );
  OR2V2_8TH40 U21 ( .A1(carry[21]), .A2(A[21]), .Z(carry[22]) );
  OR2V2_8TH40 U22 ( .A1(carry[23]), .A2(A[23]), .Z(carry[24]) );
  OR2V2_8TH40 U23 ( .A1(carry[24]), .A2(A[24]), .Z(carry[25]) );
  OR2V2_8TH40 U24 ( .A1(carry[25]), .A2(A[25]), .Z(carry[26]) );
  OR2V2_8TH40 U25 ( .A1(carry[28]), .A2(A[28]), .Z(carry[29]) );
  OR2V2_8TH40 U26 ( .A1(carry[15]), .A2(A[15]), .Z(carry[16]) );
  OR2V2_8TH40 U27 ( .A1(carry[22]), .A2(A[22]), .Z(carry[23]) );
  OR2V2_8TH40 U28 ( .A1(carry[26]), .A2(A[26]), .Z(carry[27]) );
  OR2V2_8TH40 U29 ( .A1(carry[27]), .A2(A[27]), .Z(carry[28]) );
  OR2V2_8TH40 U30 ( .A1(carry[29]), .A2(A[29]), .Z(carry[30]) );
  OR2V2_8TH40 U31 ( .A1(A[2]), .A2(n3), .Z(carry[3]) );
  INV2_8TH40 U32 ( .I(B[2]), .ZN(n3) );
  XNOR2V2_8TH40 U33 ( .A1(carry[10]), .A2(A[10]), .ZN(DIFF[10]) );
  XNOR2V2_8TH40 U34 ( .A1(carry[11]), .A2(A[11]), .ZN(DIFF[11]) );
  XNOR2V2_8TH40 U35 ( .A1(carry[12]), .A2(A[12]), .ZN(DIFF[12]) );
  XNOR2V2_8TH40 U36 ( .A1(carry[13]), .A2(A[13]), .ZN(DIFF[13]) );
  XNOR2V2_8TH40 U37 ( .A1(carry[14]), .A2(A[14]), .ZN(DIFF[14]) );
  XNOR2V2_8TH40 U38 ( .A1(carry[15]), .A2(A[15]), .ZN(DIFF[15]) );
  XNOR2V2_8TH40 U39 ( .A1(carry[16]), .A2(A[16]), .ZN(DIFF[16]) );
  XNOR2V2_8TH40 U40 ( .A1(carry[17]), .A2(A[17]), .ZN(DIFF[17]) );
  XNOR2V2_8TH40 U41 ( .A1(carry[18]), .A2(A[18]), .ZN(DIFF[18]) );
  XNOR2V2_8TH40 U42 ( .A1(carry[19]), .A2(A[19]), .ZN(DIFF[19]) );
  XNOR2V2_8TH40 U43 ( .A1(carry[20]), .A2(A[20]), .ZN(DIFF[20]) );
  XNOR2V2_8TH40 U44 ( .A1(carry[21]), .A2(A[21]), .ZN(DIFF[21]) );
  XNOR2V2_8TH40 U45 ( .A1(carry[22]), .A2(A[22]), .ZN(DIFF[22]) );
  XNOR2V2_8TH40 U46 ( .A1(carry[23]), .A2(A[23]), .ZN(DIFF[23]) );
  XNOR2V2_8TH40 U47 ( .A1(carry[24]), .A2(A[24]), .ZN(DIFF[24]) );
  XNOR2V2_8TH40 U48 ( .A1(carry[25]), .A2(A[25]), .ZN(DIFF[25]) );
  XNOR2V2_8TH40 U49 ( .A1(carry[26]), .A2(A[26]), .ZN(DIFF[26]) );
  XNOR2V2_8TH40 U50 ( .A1(carry[27]), .A2(A[27]), .ZN(DIFF[27]) );
  XNOR2V2_8TH40 U51 ( .A1(carry[28]), .A2(A[28]), .ZN(DIFF[28]) );
  XNOR2V2_8TH40 U52 ( .A1(carry[29]), .A2(A[29]), .ZN(DIFF[29]) );
  XNOR2V2_8TH40 U53 ( .A1(carry[30]), .A2(A[30]), .ZN(DIFF[30]) );
  XNOR2V2_8TH40 U54 ( .A1(A[31]), .A2(carry[31]), .ZN(DIFF[31]) );
  XNOR2V2_8TH40 U55 ( .A1(carry[3]), .A2(A[3]), .ZN(DIFF[3]) );
  XNOR2V2_8TH40 U56 ( .A1(carry[4]), .A2(A[4]), .ZN(DIFF[4]) );
  XNOR2V2_8TH40 U57 ( .A1(carry[5]), .A2(A[5]), .ZN(DIFF[5]) );
  XNOR2V2_8TH40 U58 ( .A1(carry[6]), .A2(A[6]), .ZN(DIFF[6]) );
  XNOR2V2_8TH40 U59 ( .A1(carry[7]), .A2(A[7]), .ZN(DIFF[7]) );
  XNOR2V2_8TH40 U60 ( .A1(carry[8]), .A2(A[8]), .ZN(DIFF[8]) );
  XNOR2V2_8TH40 U61 ( .A1(carry[9]), .A2(A[9]), .ZN(DIFF[9]) );
  XNOR2V2_8TH40 U62 ( .A1(A[2]), .A2(n3), .ZN(DIFF[2]) );
endmodule


module coprocessor0 ( clk, rst, cp0_reg_we, cp0_reg_waddr, cp0_reg_raddr, 
        cp0_reg_wdata, int_i, except_type_i, cur_inst_addr_i, in_delayslot_i, 
        cp0_reg_rdata, count_reg, compare_reg, status_reg, cause_reg, epc_reg, 
        config_reg, prid_reg, timer_int_o );
  input [4:0] cp0_reg_waddr;
  input [4:0] cp0_reg_raddr;
  input [31:0] cp0_reg_wdata;
  input [5:0] int_i;
  input [31:0] except_type_i;
  input [31:0] cur_inst_addr_i;
  output [31:0] cp0_reg_rdata;
  output [31:0] count_reg;
  output [31:0] compare_reg;
  output [31:0] status_reg;
  output [31:0] cause_reg;
  output [31:0] epc_reg;
  output [31:0] config_reg;
  output [31:0] prid_reg;
  input clk, rst, cp0_reg_we, in_delayslot_i;
  output timer_int_o;
  wire   N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N290, N291, N292, N293, N294, N295, N296,
         N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307,
         N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318,
         N319, N320, N321, N683, N684, N685, N686, N687, N688, N689, N690,
         N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701,
         N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, N712,
         N713, N714, N867, N868, N869, N870, N871, N872, N873, N874, N875,
         N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886,
         N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897,
         N898, N899, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225;

  DQV4_8TH40 count_reg_reg_0_ ( .D(N683), .CK(clk), .Q(count_reg[0]) );
  DQV4_8TH40 count_reg_reg_1_ ( .D(N684), .CK(clk), .Q(count_reg[1]) );
  DQV4_8TH40 count_reg_reg_2_ ( .D(N685), .CK(clk), .Q(count_reg[2]) );
  DQV4_8TH40 count_reg_reg_3_ ( .D(N686), .CK(clk), .Q(count_reg[3]) );
  DQV4_8TH40 count_reg_reg_4_ ( .D(N687), .CK(clk), .Q(count_reg[4]) );
  DQV4_8TH40 count_reg_reg_5_ ( .D(N688), .CK(clk), .Q(count_reg[5]) );
  DQV4_8TH40 count_reg_reg_6_ ( .D(N689), .CK(clk), .Q(count_reg[6]) );
  DQV4_8TH40 count_reg_reg_7_ ( .D(N690), .CK(clk), .Q(count_reg[7]) );
  DQV4_8TH40 count_reg_reg_8_ ( .D(N691), .CK(clk), .Q(count_reg[8]) );
  DQV4_8TH40 count_reg_reg_9_ ( .D(N692), .CK(clk), .Q(count_reg[9]) );
  DQV4_8TH40 count_reg_reg_10_ ( .D(N693), .CK(clk), .Q(count_reg[10]) );
  DQV4_8TH40 count_reg_reg_11_ ( .D(N694), .CK(clk), .Q(count_reg[11]) );
  DQV4_8TH40 count_reg_reg_12_ ( .D(N695), .CK(clk), .Q(count_reg[12]) );
  DQV4_8TH40 count_reg_reg_13_ ( .D(N696), .CK(clk), .Q(count_reg[13]) );
  DQV4_8TH40 count_reg_reg_14_ ( .D(N697), .CK(clk), .Q(count_reg[14]) );
  DQV4_8TH40 count_reg_reg_15_ ( .D(N698), .CK(clk), .Q(count_reg[15]) );
  DQV4_8TH40 count_reg_reg_16_ ( .D(N699), .CK(clk), .Q(count_reg[16]) );
  DQV4_8TH40 count_reg_reg_17_ ( .D(N700), .CK(clk), .Q(count_reg[17]) );
  DQV4_8TH40 count_reg_reg_18_ ( .D(N701), .CK(clk), .Q(count_reg[18]) );
  DQV4_8TH40 count_reg_reg_19_ ( .D(N702), .CK(clk), .Q(count_reg[19]) );
  DQV4_8TH40 count_reg_reg_20_ ( .D(N703), .CK(clk), .Q(count_reg[20]) );
  DQV4_8TH40 count_reg_reg_21_ ( .D(N704), .CK(clk), .Q(count_reg[21]) );
  DQV4_8TH40 count_reg_reg_22_ ( .D(N705), .CK(clk), .Q(count_reg[22]) );
  DQV4_8TH40 count_reg_reg_23_ ( .D(N706), .CK(clk), .Q(count_reg[23]) );
  DQV4_8TH40 count_reg_reg_24_ ( .D(N707), .CK(clk), .Q(count_reg[24]) );
  DQV4_8TH40 count_reg_reg_25_ ( .D(N708), .CK(clk), .Q(count_reg[25]) );
  DQV4_8TH40 count_reg_reg_26_ ( .D(N709), .CK(clk), .Q(count_reg[26]) );
  DQV4_8TH40 count_reg_reg_27_ ( .D(N710), .CK(clk), .Q(count_reg[27]) );
  DQV4_8TH40 count_reg_reg_28_ ( .D(N711), .CK(clk), .Q(count_reg[28]) );
  DQV4_8TH40 count_reg_reg_29_ ( .D(N712), .CK(clk), .Q(count_reg[29]) );
  DQV4_8TH40 count_reg_reg_30_ ( .D(N713), .CK(clk), .Q(count_reg[30]) );
  DQV4_8TH40 count_reg_reg_31_ ( .D(N714), .CK(clk), .Q(count_reg[31]) );
  DQV4_8TH40 cause_reg_reg_5_ ( .D(n395), .CK(clk), .Q(cause_reg[5]) );
  DQV4_8TH40 cause_reg_reg_4_ ( .D(n396), .CK(clk), .Q(cause_reg[4]) );
  DQV4_8TH40 cause_reg_reg_3_ ( .D(n397), .CK(clk), .Q(cause_reg[3]) );
  DQV4_8TH40 cause_reg_reg_2_ ( .D(n398), .CK(clk), .Q(cause_reg[2]) );
  DQV4_8TH40 compare_reg_reg_31_ ( .D(n462), .CK(clk), .Q(compare_reg[31]) );
  DQV4_8TH40 compare_reg_reg_30_ ( .D(n461), .CK(clk), .Q(compare_reg[30]) );
  DQV4_8TH40 compare_reg_reg_29_ ( .D(n460), .CK(clk), .Q(compare_reg[29]) );
  DQV4_8TH40 compare_reg_reg_28_ ( .D(n459), .CK(clk), .Q(compare_reg[28]) );
  DQV4_8TH40 compare_reg_reg_27_ ( .D(n458), .CK(clk), .Q(compare_reg[27]) );
  DQV4_8TH40 compare_reg_reg_26_ ( .D(n457), .CK(clk), .Q(compare_reg[26]) );
  DQV4_8TH40 compare_reg_reg_25_ ( .D(n456), .CK(clk), .Q(compare_reg[25]) );
  DQV4_8TH40 compare_reg_reg_24_ ( .D(n455), .CK(clk), .Q(compare_reg[24]) );
  DQV4_8TH40 compare_reg_reg_23_ ( .D(n454), .CK(clk), .Q(compare_reg[23]) );
  DQV4_8TH40 compare_reg_reg_22_ ( .D(n453), .CK(clk), .Q(compare_reg[22]) );
  DQV4_8TH40 compare_reg_reg_21_ ( .D(n452), .CK(clk), .Q(compare_reg[21]) );
  DQV4_8TH40 compare_reg_reg_20_ ( .D(n451), .CK(clk), .Q(compare_reg[20]) );
  DQV4_8TH40 compare_reg_reg_19_ ( .D(n450), .CK(clk), .Q(compare_reg[19]) );
  DQV4_8TH40 compare_reg_reg_18_ ( .D(n449), .CK(clk), .Q(compare_reg[18]) );
  DQV4_8TH40 compare_reg_reg_17_ ( .D(n448), .CK(clk), .Q(compare_reg[17]) );
  DQV4_8TH40 compare_reg_reg_16_ ( .D(n447), .CK(clk), .Q(compare_reg[16]) );
  DQV4_8TH40 compare_reg_reg_15_ ( .D(n446), .CK(clk), .Q(compare_reg[15]) );
  DQV4_8TH40 compare_reg_reg_14_ ( .D(n445), .CK(clk), .Q(compare_reg[14]) );
  DQV4_8TH40 compare_reg_reg_13_ ( .D(n444), .CK(clk), .Q(compare_reg[13]) );
  DQV4_8TH40 compare_reg_reg_12_ ( .D(n443), .CK(clk), .Q(compare_reg[12]) );
  DQV4_8TH40 compare_reg_reg_11_ ( .D(n442), .CK(clk), .Q(compare_reg[11]) );
  DQV4_8TH40 compare_reg_reg_10_ ( .D(n441), .CK(clk), .Q(compare_reg[10]) );
  DQV4_8TH40 compare_reg_reg_9_ ( .D(n440), .CK(clk), .Q(compare_reg[9]) );
  DQV4_8TH40 compare_reg_reg_8_ ( .D(n439), .CK(clk), .Q(compare_reg[8]) );
  DQV4_8TH40 compare_reg_reg_7_ ( .D(n438), .CK(clk), .Q(compare_reg[7]) );
  DQV4_8TH40 compare_reg_reg_6_ ( .D(n437), .CK(clk), .Q(compare_reg[6]) );
  DQV4_8TH40 compare_reg_reg_5_ ( .D(n436), .CK(clk), .Q(compare_reg[5]) );
  DQV4_8TH40 compare_reg_reg_4_ ( .D(n435), .CK(clk), .Q(compare_reg[4]) );
  DQV4_8TH40 compare_reg_reg_3_ ( .D(n434), .CK(clk), .Q(compare_reg[3]) );
  DQV4_8TH40 compare_reg_reg_2_ ( .D(n433), .CK(clk), .Q(compare_reg[2]) );
  DQV4_8TH40 compare_reg_reg_1_ ( .D(n432), .CK(clk), .Q(compare_reg[1]) );
  DQV4_8TH40 compare_reg_reg_0_ ( .D(n431), .CK(clk), .Q(compare_reg[0]) );
  DQV4_8TH40 timer_int_o_reg ( .D(n430), .CK(clk), .Q(timer_int_o) );
  DQV4_8TH40 status_reg_reg_31_ ( .D(n429), .CK(clk), .Q(status_reg[31]) );
  DQV4_8TH40 status_reg_reg_30_ ( .D(n428), .CK(clk), .Q(status_reg[30]) );
  DQV4_8TH40 status_reg_reg_29_ ( .D(n427), .CK(clk), .Q(status_reg[29]) );
  DQV4_8TH40 status_reg_reg_28_ ( .D(n426), .CK(clk), .Q(status_reg[28]) );
  DQV4_8TH40 status_reg_reg_27_ ( .D(n425), .CK(clk), .Q(status_reg[27]) );
  DQV4_8TH40 status_reg_reg_26_ ( .D(n424), .CK(clk), .Q(status_reg[26]) );
  DQV4_8TH40 status_reg_reg_25_ ( .D(n423), .CK(clk), .Q(status_reg[25]) );
  DQV4_8TH40 status_reg_reg_24_ ( .D(n422), .CK(clk), .Q(status_reg[24]) );
  DQV4_8TH40 status_reg_reg_23_ ( .D(n421), .CK(clk), .Q(status_reg[23]) );
  DQV4_8TH40 status_reg_reg_22_ ( .D(n420), .CK(clk), .Q(status_reg[22]) );
  DQV4_8TH40 status_reg_reg_21_ ( .D(n419), .CK(clk), .Q(status_reg[21]) );
  DQV4_8TH40 status_reg_reg_20_ ( .D(n418), .CK(clk), .Q(status_reg[20]) );
  DQV4_8TH40 status_reg_reg_19_ ( .D(n417), .CK(clk), .Q(status_reg[19]) );
  DQV4_8TH40 status_reg_reg_18_ ( .D(n416), .CK(clk), .Q(status_reg[18]) );
  DQV4_8TH40 status_reg_reg_17_ ( .D(n415), .CK(clk), .Q(status_reg[17]) );
  DQV4_8TH40 status_reg_reg_16_ ( .D(n414), .CK(clk), .Q(status_reg[16]) );
  DQV4_8TH40 status_reg_reg_15_ ( .D(n413), .CK(clk), .Q(status_reg[15]) );
  DQV4_8TH40 status_reg_reg_14_ ( .D(n412), .CK(clk), .Q(status_reg[14]) );
  DQV4_8TH40 status_reg_reg_13_ ( .D(n411), .CK(clk), .Q(status_reg[13]) );
  DQV4_8TH40 status_reg_reg_12_ ( .D(n410), .CK(clk), .Q(status_reg[12]) );
  DQV4_8TH40 status_reg_reg_11_ ( .D(n409), .CK(clk), .Q(status_reg[11]) );
  DQV4_8TH40 status_reg_reg_10_ ( .D(n408), .CK(clk), .Q(status_reg[10]) );
  DQV4_8TH40 status_reg_reg_9_ ( .D(n407), .CK(clk), .Q(status_reg[9]) );
  DQV4_8TH40 status_reg_reg_8_ ( .D(n406), .CK(clk), .Q(status_reg[8]) );
  DQV4_8TH40 status_reg_reg_7_ ( .D(n405), .CK(clk), .Q(status_reg[7]) );
  DQV4_8TH40 status_reg_reg_6_ ( .D(n404), .CK(clk), .Q(status_reg[6]) );
  DQV4_8TH40 status_reg_reg_5_ ( .D(n403), .CK(clk), .Q(status_reg[5]) );
  DQV4_8TH40 status_reg_reg_4_ ( .D(n402), .CK(clk), .Q(status_reg[4]) );
  DQV4_8TH40 status_reg_reg_3_ ( .D(n401), .CK(clk), .Q(status_reg[3]) );
  DQV4_8TH40 status_reg_reg_2_ ( .D(n400), .CK(clk), .Q(status_reg[2]) );
  DQV4_8TH40 status_reg_reg_1_ ( .D(n399), .CK(clk), .Q(status_reg[1]) );
  DQV4_8TH40 epc_reg_reg_31_ ( .D(n362), .CK(clk), .Q(epc_reg[31]) );
  DQV4_8TH40 epc_reg_reg_30_ ( .D(n363), .CK(clk), .Q(epc_reg[30]) );
  DQV4_8TH40 epc_reg_reg_29_ ( .D(n364), .CK(clk), .Q(epc_reg[29]) );
  DQV4_8TH40 epc_reg_reg_28_ ( .D(n365), .CK(clk), .Q(epc_reg[28]) );
  DQV4_8TH40 epc_reg_reg_27_ ( .D(n366), .CK(clk), .Q(epc_reg[27]) );
  DQV4_8TH40 epc_reg_reg_26_ ( .D(n367), .CK(clk), .Q(epc_reg[26]) );
  DQV4_8TH40 epc_reg_reg_25_ ( .D(n368), .CK(clk), .Q(epc_reg[25]) );
  DQV4_8TH40 epc_reg_reg_24_ ( .D(n369), .CK(clk), .Q(epc_reg[24]) );
  DQV4_8TH40 epc_reg_reg_23_ ( .D(n370), .CK(clk), .Q(epc_reg[23]) );
  DQV4_8TH40 epc_reg_reg_22_ ( .D(n371), .CK(clk), .Q(epc_reg[22]) );
  DQV4_8TH40 epc_reg_reg_21_ ( .D(n372), .CK(clk), .Q(epc_reg[21]) );
  DQV4_8TH40 epc_reg_reg_20_ ( .D(n373), .CK(clk), .Q(epc_reg[20]) );
  DQV4_8TH40 epc_reg_reg_19_ ( .D(n374), .CK(clk), .Q(epc_reg[19]) );
  DQV4_8TH40 epc_reg_reg_18_ ( .D(n375), .CK(clk), .Q(epc_reg[18]) );
  DQV4_8TH40 epc_reg_reg_17_ ( .D(n376), .CK(clk), .Q(epc_reg[17]) );
  DQV4_8TH40 epc_reg_reg_16_ ( .D(n377), .CK(clk), .Q(epc_reg[16]) );
  DQV4_8TH40 epc_reg_reg_15_ ( .D(n378), .CK(clk), .Q(epc_reg[15]) );
  DQV4_8TH40 epc_reg_reg_14_ ( .D(n379), .CK(clk), .Q(epc_reg[14]) );
  DQV4_8TH40 epc_reg_reg_13_ ( .D(n380), .CK(clk), .Q(epc_reg[13]) );
  DQV4_8TH40 epc_reg_reg_12_ ( .D(n381), .CK(clk), .Q(epc_reg[12]) );
  DQV4_8TH40 epc_reg_reg_11_ ( .D(n382), .CK(clk), .Q(epc_reg[11]) );
  DQV4_8TH40 epc_reg_reg_10_ ( .D(n383), .CK(clk), .Q(epc_reg[10]) );
  DQV4_8TH40 epc_reg_reg_9_ ( .D(n384), .CK(clk), .Q(epc_reg[9]) );
  DQV4_8TH40 epc_reg_reg_8_ ( .D(n385), .CK(clk), .Q(epc_reg[8]) );
  DQV4_8TH40 epc_reg_reg_7_ ( .D(n386), .CK(clk), .Q(epc_reg[7]) );
  DQV4_8TH40 epc_reg_reg_6_ ( .D(n387), .CK(clk), .Q(epc_reg[6]) );
  DQV4_8TH40 epc_reg_reg_5_ ( .D(n388), .CK(clk), .Q(epc_reg[5]) );
  DQV4_8TH40 epc_reg_reg_4_ ( .D(n389), .CK(clk), .Q(epc_reg[4]) );
  DQV4_8TH40 epc_reg_reg_3_ ( .D(n390), .CK(clk), .Q(epc_reg[3]) );
  DQV4_8TH40 epc_reg_reg_2_ ( .D(n391), .CK(clk), .Q(epc_reg[2]) );
  DQV4_8TH40 epc_reg_reg_1_ ( .D(n392), .CK(clk), .Q(epc_reg[1]) );
  DQV4_8TH40 epc_reg_reg_0_ ( .D(n393), .CK(clk), .Q(epc_reg[0]) );
  DQV4_8TH40 cause_reg_reg_31_ ( .D(n394), .CK(clk), .Q(cause_reg[31]) );
  DQV4_8TH40 status_reg_reg_0_ ( .D(n361), .CK(clk), .Q(status_reg[0]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_31_ ( .E(N867), .D(N899), .Q(
        cp0_reg_rdata[31]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_30_ ( .E(N867), .D(N898), .Q(
        cp0_reg_rdata[30]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_28_ ( .E(N867), .D(N896), .Q(
        cp0_reg_rdata[28]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_23_ ( .E(N867), .D(N891), .Q(
        cp0_reg_rdata[23]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_21_ ( .E(N867), .D(N889), .Q(
        cp0_reg_rdata[21]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_19_ ( .E(N867), .D(N887), .Q(
        cp0_reg_rdata[19]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_18_ ( .E(N867), .D(N886), .Q(
        cp0_reg_rdata[18]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_17_ ( .E(N867), .D(N885), .Q(
        cp0_reg_rdata[17]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_16_ ( .E(N867), .D(N884), .Q(
        cp0_reg_rdata[16]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_15_ ( .E(N867), .D(N883), .Q(
        cp0_reg_rdata[15]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_14_ ( .E(N867), .D(N882), .Q(
        cp0_reg_rdata[14]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_13_ ( .E(N867), .D(N881), .Q(
        cp0_reg_rdata[13]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_12_ ( .E(N867), .D(N880), .Q(
        cp0_reg_rdata[12]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_11_ ( .E(N867), .D(N879), .Q(
        cp0_reg_rdata[11]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_10_ ( .E(N867), .D(N878), .Q(
        cp0_reg_rdata[10]) );
  LAHQV1_8TH40 cp0_reg_rdata_reg_9_ ( .E(N867), .D(N877), .Q(cp0_reg_rdata[9])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_8_ ( .E(N867), .D(N876), .Q(cp0_reg_rdata[8])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_7_ ( .E(N867), .D(N875), .Q(cp0_reg_rdata[7])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_6_ ( .E(N867), .D(N874), .Q(cp0_reg_rdata[6])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_4_ ( .E(N867), .D(N872), .Q(cp0_reg_rdata[4])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_3_ ( .E(N867), .D(N871), .Q(cp0_reg_rdata[3])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_2_ ( .E(N867), .D(N870), .Q(cp0_reg_rdata[2])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_1_ ( .E(N867), .D(N869), .Q(cp0_reg_rdata[1])
         );
  LAHQV1_8TH40 cp0_reg_rdata_reg_0_ ( .E(N867), .D(N868), .Q(cp0_reg_rdata[0])
         );
  coprocessor0_DW01_cmp6_0 eq_51 ( .A(count_reg), .B(compare_reg), .TC(1'b0), 
        .EQ(N62) );
  coprocessor0_DW01_inc_0 add_48 ( .A(count_reg), .SUM({N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30})
         );
  coprocessor0_DW01_sub_0 r123 ( .A(cur_inst_addr_i), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, in_delayslot_i, 1'b0, 1'b0}), .CI(1'b0), .DIFF({N321, N320, 
        N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, 
        N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290}) );
  EDGRNQV2_8TH40 cause_reg_reg_23_ ( .RN(n225), .D(cp0_reg_wdata[23]), .E(n224), .CK(clk), .Q(cause_reg[23]) );
  EDGRNQV2_8TH40 cause_reg_reg_22_ ( .RN(n225), .D(cp0_reg_wdata[22]), .E(n224), .CK(clk), .Q(cause_reg[22]) );
  EDGRNQV2_8TH40 cause_reg_reg_9_ ( .RN(n225), .D(cp0_reg_wdata[9]), .E(n224), 
        .CK(clk), .Q(cause_reg[9]) );
  EDGRNQV2_8TH40 cause_reg_reg_8_ ( .RN(n225), .D(cp0_reg_wdata[8]), .E(n224), 
        .CK(clk), .Q(cause_reg[8]) );
  DGRNQV2_8TH40 cause_reg_reg_15_ ( .D(int_i[5]), .RN(n225), .CK(clk), .Q(
        cause_reg[15]) );
  DGRNQV2_8TH40 cause_reg_reg_14_ ( .D(int_i[4]), .RN(n225), .CK(clk), .Q(
        cause_reg[14]) );
  DGRNQV2_8TH40 cause_reg_reg_13_ ( .D(int_i[3]), .RN(n225), .CK(clk), .Q(
        cause_reg[13]) );
  DGRNQV2_8TH40 cause_reg_reg_12_ ( .D(int_i[2]), .RN(n225), .CK(clk), .Q(
        cause_reg[12]) );
  DGRNQV2_8TH40 cause_reg_reg_11_ ( .D(int_i[1]), .RN(n225), .CK(clk), .Q(
        cause_reg[11]) );
  DGRNQV2_8TH40 cause_reg_reg_10_ ( .D(int_i[0]), .RN(n225), .CK(clk), .Q(
        cause_reg[10]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_29_ ( .E(N867), .D(N897), .Q(
        cp0_reg_rdata[29]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_27_ ( .E(N867), .D(N895), .Q(
        cp0_reg_rdata[27]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_26_ ( .E(N867), .D(N894), .Q(
        cp0_reg_rdata[26]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_25_ ( .E(N867), .D(N893), .Q(
        cp0_reg_rdata[25]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_24_ ( .E(N867), .D(N892), .Q(
        cp0_reg_rdata[24]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_22_ ( .E(N867), .D(N890), .Q(
        cp0_reg_rdata[22]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_20_ ( .E(N867), .D(N888), .Q(
        cp0_reg_rdata[20]) );
  LAHQV4_8TH40 cp0_reg_rdata_reg_5_ ( .E(N867), .D(N873), .Q(cp0_reg_rdata[5])
         );
  AO222V4_8TH40 U3 ( .A1(N292), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[2]), 
        .C1(epc_reg[2]), .C2(n139), .Z(n391) );
  AO222V4_8TH40 U4 ( .A1(N293), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[3]), 
        .C1(epc_reg[3]), .C2(n139), .Z(n390) );
  AO222V4_8TH40 U5 ( .A1(N294), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[4]), 
        .C1(epc_reg[4]), .C2(n139), .Z(n389) );
  AO222V4_8TH40 U6 ( .A1(N295), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[5]), 
        .C1(epc_reg[5]), .C2(n139), .Z(n388) );
  AO222V4_8TH40 U7 ( .A1(N296), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[6]), 
        .C1(epc_reg[6]), .C2(n139), .Z(n387) );
  AO222V4_8TH40 U8 ( .A1(N297), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[7]), 
        .C1(epc_reg[7]), .C2(n139), .Z(n386) );
  AO222V4_8TH40 U9 ( .A1(N298), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[8]), 
        .C1(epc_reg[8]), .C2(n139), .Z(n385) );
  AO222V4_8TH40 U10 ( .A1(N299), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[9]), 
        .C1(epc_reg[9]), .C2(n139), .Z(n384) );
  AO222V4_8TH40 U11 ( .A1(N300), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[10]), 
        .C1(epc_reg[10]), .C2(n139), .Z(n383) );
  AO222V4_8TH40 U14 ( .A1(N301), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[11]), 
        .C1(epc_reg[11]), .C2(n139), .Z(n382) );
  AO222V4_8TH40 U15 ( .A1(N302), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[12]), 
        .C1(epc_reg[12]), .C2(n139), .Z(n381) );
  AO222V4_8TH40 U16 ( .A1(N303), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[13]), 
        .C1(epc_reg[13]), .C2(n139), .Z(n380) );
  AO222V4_8TH40 U17 ( .A1(N304), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[14]), 
        .C1(epc_reg[14]), .C2(n139), .Z(n379) );
  AO222V4_8TH40 U18 ( .A1(N305), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[15]), 
        .C1(epc_reg[15]), .C2(n139), .Z(n378) );
  AO222V4_8TH40 U19 ( .A1(N306), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[16]), 
        .C1(epc_reg[16]), .C2(n139), .Z(n377) );
  AO222V4_8TH40 U20 ( .A1(N307), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[17]), 
        .C1(epc_reg[17]), .C2(n139), .Z(n376) );
  AO222V4_8TH40 U21 ( .A1(N308), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[18]), 
        .C1(epc_reg[18]), .C2(n139), .Z(n375) );
  AO222V4_8TH40 U22 ( .A1(N309), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[19]), 
        .C1(epc_reg[19]), .C2(n139), .Z(n374) );
  AO222V4_8TH40 U23 ( .A1(N310), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[20]), 
        .C1(epc_reg[20]), .C2(n139), .Z(n373) );
  AO222V4_8TH40 U24 ( .A1(N311), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[21]), 
        .C1(epc_reg[21]), .C2(n139), .Z(n372) );
  AO222V4_8TH40 U25 ( .A1(N312), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[22]), 
        .C1(epc_reg[22]), .C2(n139), .Z(n371) );
  AO222V4_8TH40 U26 ( .A1(N313), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[23]), 
        .C1(epc_reg[23]), .C2(n139), .Z(n370) );
  AO222V4_8TH40 U27 ( .A1(N314), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[24]), 
        .C1(epc_reg[24]), .C2(n139), .Z(n369) );
  AO222V4_8TH40 U28 ( .A1(N315), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[25]), 
        .C1(epc_reg[25]), .C2(n139), .Z(n368) );
  AO222V4_8TH40 U29 ( .A1(N316), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[26]), 
        .C1(epc_reg[26]), .C2(n139), .Z(n367) );
  AO222V4_8TH40 U30 ( .A1(N317), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[27]), 
        .C1(epc_reg[27]), .C2(n139), .Z(n366) );
  AO222V4_8TH40 U31 ( .A1(N318), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[28]), 
        .C1(epc_reg[28]), .C2(n139), .Z(n365) );
  AO222V4_8TH40 U32 ( .A1(N319), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[29]), 
        .C1(epc_reg[29]), .C2(n139), .Z(n364) );
  AO222V4_8TH40 U33 ( .A1(N320), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[30]), 
        .C1(epc_reg[30]), .C2(n139), .Z(n363) );
  AO222V4_8TH40 U34 ( .A1(N321), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[31]), 
        .C1(epc_reg[31]), .C2(n139), .Z(n362) );
  MOAI22V4_8TH40 U35 ( .A1(n9), .A2(n221), .B1(N60), .B2(n222), .ZN(N713) );
  MOAI22V4_8TH40 U36 ( .A1(n11), .A2(n221), .B1(N59), .B2(n222), .ZN(N712) );
  MOAI22V4_8TH40 U37 ( .A1(n13), .A2(n221), .B1(N58), .B2(n222), .ZN(N711) );
  MOAI22V4_8TH40 U38 ( .A1(n15), .A2(n221), .B1(N57), .B2(n222), .ZN(N710) );
  MOAI22V4_8TH40 U39 ( .A1(n17), .A2(n221), .B1(N56), .B2(n222), .ZN(N709) );
  MOAI22V4_8TH40 U40 ( .A1(n19), .A2(n221), .B1(N55), .B2(n222), .ZN(N708) );
  MOAI22V4_8TH40 U41 ( .A1(n21), .A2(n221), .B1(N54), .B2(n222), .ZN(N707) );
  MOAI22V4_8TH40 U42 ( .A1(n23), .A2(n221), .B1(N53), .B2(n222), .ZN(N706) );
  MOAI22V4_8TH40 U43 ( .A1(n25), .A2(n221), .B1(N52), .B2(n222), .ZN(N705) );
  MOAI22V4_8TH40 U44 ( .A1(n27), .A2(n221), .B1(N51), .B2(n222), .ZN(N704) );
  MOAI22V4_8TH40 U45 ( .A1(n29), .A2(n221), .B1(N50), .B2(n222), .ZN(N703) );
  MOAI22V4_8TH40 U46 ( .A1(n31), .A2(n221), .B1(N49), .B2(n222), .ZN(N702) );
  MOAI22V4_8TH40 U47 ( .A1(n33), .A2(n221), .B1(N48), .B2(n222), .ZN(N701) );
  MOAI22V4_8TH40 U48 ( .A1(n35), .A2(n221), .B1(N47), .B2(n222), .ZN(N700) );
  MOAI22V4_8TH40 U49 ( .A1(n37), .A2(n221), .B1(N46), .B2(n222), .ZN(N699) );
  MOAI22V4_8TH40 U50 ( .A1(n39), .A2(n221), .B1(N45), .B2(n222), .ZN(N698) );
  MOAI22V4_8TH40 U51 ( .A1(n41), .A2(n221), .B1(N44), .B2(n222), .ZN(N697) );
  MOAI22V4_8TH40 U52 ( .A1(n43), .A2(n221), .B1(N43), .B2(n222), .ZN(N696) );
  MOAI22V4_8TH40 U53 ( .A1(n45), .A2(n221), .B1(N42), .B2(n222), .ZN(N695) );
  MOAI22V4_8TH40 U54 ( .A1(n47), .A2(n221), .B1(N41), .B2(n222), .ZN(N694) );
  MOAI22V4_8TH40 U55 ( .A1(n49), .A2(n221), .B1(N40), .B2(n222), .ZN(N693) );
  MOAI22V4_8TH40 U56 ( .A1(n51), .A2(n221), .B1(N39), .B2(n222), .ZN(N692) );
  MOAI22V4_8TH40 U57 ( .A1(n53), .A2(n221), .B1(N38), .B2(n222), .ZN(N691) );
  MOAI22V4_8TH40 U58 ( .A1(n55), .A2(n221), .B1(N37), .B2(n222), .ZN(N690) );
  MOAI22V4_8TH40 U59 ( .A1(n57), .A2(n221), .B1(N36), .B2(n222), .ZN(N689) );
  MOAI22V4_8TH40 U60 ( .A1(n59), .A2(n221), .B1(N35), .B2(n222), .ZN(N688) );
  MOAI22V4_8TH40 U61 ( .A1(n61), .A2(n221), .B1(N34), .B2(n222), .ZN(N687) );
  MOAI22V4_8TH40 U62 ( .A1(n63), .A2(n221), .B1(N33), .B2(n222), .ZN(N686) );
  MOAI22V4_8TH40 U63 ( .A1(n65), .A2(n221), .B1(N32), .B2(n222), .ZN(N685) );
  MOAI22V4_8TH40 U64 ( .A1(n67), .A2(n221), .B1(N31), .B2(n222), .ZN(N684) );
  MOAI22V4_8TH40 U65 ( .A1(n7), .A2(n221), .B1(N61), .B2(n222), .ZN(N714) );
  MOAI22V4_8TH40 U66 ( .A1(n69), .A2(n221), .B1(N30), .B2(n222), .ZN(N683) );
  MUX2NV2_8TH40 U67 ( .I0(n4), .I1(n70), .S(n71), .ZN(n430) );
  MUX2NV2_8TH40 U68 ( .I0(n89), .I1(n90), .S(n84), .ZN(n426) );
  MUX2NV2_8TH40 U69 ( .I0(n117), .I1(n118), .S(n119), .ZN(n399) );
  AOI21V2_8TH40 U70 ( .A1(except_type_i[0]), .A2(except_type_i[1]), .B(n146), 
        .ZN(n125) );
  XOR2V2_8TH40 U71 ( .A1(except_type_i[3]), .A2(n147), .Z(n146) );
  NAND2V2_8TH40 U72 ( .A1(n124), .A2(n225), .ZN(n117) );
  I2NOR3V2_8TH40 U73 ( .A1(n143), .A2(n225), .B(n136), .ZN(n139) );
  NAND2V2_8TH40 U74 ( .A1(n225), .A2(n82), .ZN(n4) );
  OAI22V2_8TH40 U75 ( .A1(n84), .A2(n110), .B1(n53), .B2(n86), .ZN(n406) );
  OAI22V2_8TH40 U76 ( .A1(n84), .A2(n103), .B1(n39), .B2(n86), .ZN(n413) );
  OAI22V2_8TH40 U77 ( .A1(n84), .A2(n96), .B1(n25), .B2(n86), .ZN(n420) );
  INV2_8TH40 U78 ( .I(timer_int_o), .ZN(n70) );
  OAOI211V2_8TH40 U79 ( .A1(n72), .A2(n73), .B(N62), .C(n4), .ZN(n71) );
  NAND4V2_8TH40 U80 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(n72) );
  OAI22V2_8TH40 U81 ( .A1(n4), .A2(n68), .B1(n6), .B2(n69), .ZN(n431) );
  OAI22V2_8TH40 U82 ( .A1(n4), .A2(n64), .B1(n6), .B2(n65), .ZN(n433) );
  OAI22V2_8TH40 U83 ( .A1(n4), .A2(n62), .B1(n6), .B2(n63), .ZN(n434) );
  OAI22V2_8TH40 U84 ( .A1(n4), .A2(n60), .B1(n6), .B2(n61), .ZN(n435) );
  OAI22V2_8TH40 U85 ( .A1(n4), .A2(n58), .B1(n6), .B2(n59), .ZN(n436) );
  OAI22V2_8TH40 U86 ( .A1(n4), .A2(n52), .B1(n6), .B2(n53), .ZN(n439) );
  OAI22V2_8TH40 U87 ( .A1(n4), .A2(n50), .B1(n6), .B2(n51), .ZN(n440) );
  OAI22V2_8TH40 U88 ( .A1(n4), .A2(n48), .B1(n6), .B2(n49), .ZN(n441) );
  OAI22V2_8TH40 U89 ( .A1(n4), .A2(n46), .B1(n6), .B2(n47), .ZN(n442) );
  OAI22V2_8TH40 U90 ( .A1(n4), .A2(n44), .B1(n6), .B2(n45), .ZN(n443) );
  OAI22V2_8TH40 U91 ( .A1(n4), .A2(n42), .B1(n6), .B2(n43), .ZN(n444) );
  OAI22V2_8TH40 U92 ( .A1(n4), .A2(n40), .B1(n6), .B2(n41), .ZN(n445) );
  OAI22V2_8TH40 U93 ( .A1(n4), .A2(n32), .B1(n6), .B2(n33), .ZN(n449) );
  OAI22V2_8TH40 U94 ( .A1(n4), .A2(n24), .B1(n6), .B2(n25), .ZN(n453) );
  OAI22V2_8TH40 U95 ( .A1(n4), .A2(n22), .B1(n6), .B2(n23), .ZN(n454) );
  OAI22V2_8TH40 U96 ( .A1(n4), .A2(n20), .B1(n6), .B2(n21), .ZN(n455) );
  OAI22V2_8TH40 U97 ( .A1(n4), .A2(n5), .B1(n6), .B2(n7), .ZN(n462) );
  OAI221V2_8TH40 U98 ( .A1(n66), .A2(n156), .B1(n118), .B2(n149), .C(n212), 
        .ZN(N869) );
  OAI221V2_8TH40 U99 ( .A1(n56), .A2(n156), .B1(n112), .B2(n149), .C(n201), 
        .ZN(N874) );
  OAI221V2_8TH40 U100 ( .A1(n54), .A2(n156), .B1(n111), .B2(n149), .C(n200), 
        .ZN(N875) );
  OAI221V2_8TH40 U101 ( .A1(n36), .A2(n156), .B1(n102), .B2(n149), .C(n179), 
        .ZN(N884) );
  OAI221V2_8TH40 U102 ( .A1(n34), .A2(n156), .B1(n101), .B2(n149), .C(n178), 
        .ZN(N885) );
  OAI221V2_8TH40 U103 ( .A1(n30), .A2(n156), .B1(n99), .B2(n149), .C(n175), 
        .ZN(N887) );
  OAI221V2_8TH40 U104 ( .A1(n28), .A2(n156), .B1(n98), .B2(n149), .C(n174), 
        .ZN(N888) );
  OAI221V2_8TH40 U105 ( .A1(n26), .A2(n156), .B1(n97), .B2(n149), .C(n173), 
        .ZN(N889) );
  OAI221V2_8TH40 U106 ( .A1(n18), .A2(n156), .B1(n93), .B2(n149), .C(n162), 
        .ZN(N893) );
  OAI221V2_8TH40 U107 ( .A1(n16), .A2(n156), .B1(n92), .B2(n149), .C(n161), 
        .ZN(N894) );
  OAI221V2_8TH40 U108 ( .A1(n14), .A2(n156), .B1(n91), .B2(n149), .C(n160), 
        .ZN(N895) );
  OAI221V2_8TH40 U109 ( .A1(n12), .A2(n156), .B1(n89), .B2(n149), .C(n159), 
        .ZN(N896) );
  OAI221V2_8TH40 U110 ( .A1(n10), .A2(n156), .B1(n88), .B2(n149), .C(n158), 
        .ZN(N897) );
  OAI221V2_8TH40 U111 ( .A1(n8), .A2(n156), .B1(n87), .B2(n149), .C(n157), 
        .ZN(N898) );
  OAI211V2_8TH40 U112 ( .A1(n148), .A2(n149), .B(n213), .C(n214), .ZN(N868) );
  OAI211V2_8TH40 U113 ( .A1(n116), .A2(n149), .B(n208), .C(n209), .ZN(N870) );
  OAI211V2_8TH40 U114 ( .A1(n115), .A2(n149), .B(n206), .C(n207), .ZN(N871) );
  OAI211V2_8TH40 U115 ( .A1(n114), .A2(n149), .B(n204), .C(n205), .ZN(N872) );
  OAI211V2_8TH40 U116 ( .A1(n113), .A2(n149), .B(n202), .C(n203), .ZN(N873) );
  OAI211V2_8TH40 U117 ( .A1(n109), .A2(n149), .B(n195), .C(n196), .ZN(N877) );
  OAI211V2_8TH40 U118 ( .A1(n108), .A2(n149), .B(n193), .C(n194), .ZN(N878) );
  OAI211V2_8TH40 U119 ( .A1(n107), .A2(n149), .B(n191), .C(n192), .ZN(N879) );
  OAI211V2_8TH40 U120 ( .A1(n106), .A2(n149), .B(n189), .C(n190), .ZN(N880) );
  OAI211V2_8TH40 U121 ( .A1(n105), .A2(n149), .B(n187), .C(n188), .ZN(N881) );
  OAI211V2_8TH40 U122 ( .A1(n104), .A2(n149), .B(n185), .C(n186), .ZN(N882) );
  OAI211V2_8TH40 U123 ( .A1(n100), .A2(n149), .B(n176), .C(n177), .ZN(N886) );
  OAI211V2_8TH40 U124 ( .A1(n95), .A2(n149), .B(n166), .C(n167), .ZN(N891) );
  AOI22V2_8TH40 U125 ( .A1(cause_reg[23]), .A2(n154), .B1(n155), .B2(
        compare_reg[23]), .ZN(n166) );
  OAI211V2_8TH40 U126 ( .A1(n94), .A2(n149), .B(n163), .C(n164), .ZN(N892) );
  OAI211V2_8TH40 U127 ( .A1(n85), .A2(n149), .B(n150), .C(n151), .ZN(N899) );
  OAI211V2_8TH40 U128 ( .A1(n38), .A2(n156), .B(n180), .C(n181), .ZN(N883) );
  AOI22V2_8TH40 U129 ( .A1(n182), .A2(n183), .B1(cause_reg[15]), .B2(n154), 
        .ZN(n180) );
  OAI22V2_8TH40 U130 ( .A1(n122), .A2(n134), .B1(n127), .B2(n132), .ZN(n395)
         );
  OAI22V2_8TH40 U131 ( .A1(n122), .A2(n128), .B1(n121), .B2(n129), .ZN(n398)
         );
  OAI22V2_8TH40 U132 ( .A1(n122), .A2(n130), .B1(n131), .B2(n132), .ZN(n397)
         );
  OAI211V2_8TH40 U133 ( .A1(n197), .A2(n169), .B(n198), .C(n199), .ZN(N876) );
  OAI211V2_8TH40 U134 ( .A1(n168), .A2(n169), .B(n170), .C(n171), .ZN(N890) );
  AOI221V2_8TH40 U135 ( .A1(n155), .A2(compare_reg[22]), .B1(cause_reg[22]), 
        .B2(n154), .C(n165), .ZN(n171) );
  OAI21V2_8TH40 U136 ( .A1(n122), .A2(n133), .B(n129), .ZN(n396) );
  NAND4V2_8TH40 U137 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(n73) );
  NOR2V2_8TH40 U138 ( .A1(rst), .A2(n135), .ZN(n394) );
  INV2_8TH40 U139 ( .I(cp0_reg_raddr[3]), .ZN(n220) );
  INV2_8TH40 U140 ( .I(status_reg[6]), .ZN(n112) );
  INV2_8TH40 U141 ( .I(status_reg[7]), .ZN(n111) );
  INV2_8TH40 U142 ( .I(status_reg[16]), .ZN(n102) );
  INV2_8TH40 U143 ( .I(status_reg[17]), .ZN(n101) );
  INV2_8TH40 U144 ( .I(status_reg[19]), .ZN(n99) );
  INV2_8TH40 U145 ( .I(status_reg[20]), .ZN(n98) );
  INV2_8TH40 U146 ( .I(status_reg[21]), .ZN(n97) );
  INV2_8TH40 U147 ( .I(status_reg[25]), .ZN(n93) );
  INV2_8TH40 U148 ( .I(status_reg[26]), .ZN(n92) );
  INV2_8TH40 U149 ( .I(status_reg[27]), .ZN(n91) );
  INV2_8TH40 U150 ( .I(status_reg[29]), .ZN(n88) );
  INV2_8TH40 U151 ( .I(status_reg[30]), .ZN(n87) );
  INV2_8TH40 U152 ( .I(status_reg[18]), .ZN(n100) );
  INV2_8TH40 U153 ( .I(status_reg[24]), .ZN(n94) );
  INV2_8TH40 U154 ( .I(status_reg[2]), .ZN(n116) );
  INV2_8TH40 U155 ( .I(status_reg[3]), .ZN(n115) );
  INV2_8TH40 U156 ( .I(status_reg[4]), .ZN(n114) );
  INV2_8TH40 U157 ( .I(status_reg[5]), .ZN(n113) );
  INV2_8TH40 U158 ( .I(status_reg[23]), .ZN(n95) );
  INV2_8TH40 U159 ( .I(status_reg[31]), .ZN(n85) );
  INV2_8TH40 U160 ( .I(status_reg[28]), .ZN(n89) );
  INOR3V0_8TH40 U161 ( .A1(cp0_reg_waddr[0]), .B1(cp0_reg_waddr[1]), .B2(n3), 
        .ZN(n224) );
  CLKNV1_8TH40 U162 ( .I(compare_reg[31]), .ZN(n5) );
  OAI22V0_8TH40 U163 ( .A1(n4), .A2(n8), .B1(n6), .B2(n9), .ZN(n461) );
  OAI22V0_8TH40 U164 ( .A1(n4), .A2(n10), .B1(n6), .B2(n11), .ZN(n460) );
  OAI22V0_8TH40 U165 ( .A1(n4), .A2(n12), .B1(n6), .B2(n13), .ZN(n459) );
  OAI22V0_8TH40 U166 ( .A1(n4), .A2(n14), .B1(n6), .B2(n15), .ZN(n458) );
  OAI22V0_8TH40 U167 ( .A1(n4), .A2(n16), .B1(n6), .B2(n17), .ZN(n457) );
  OAI22V0_8TH40 U168 ( .A1(n4), .A2(n18), .B1(n6), .B2(n19), .ZN(n456) );
  CLKNV1_8TH40 U169 ( .I(compare_reg[24]), .ZN(n20) );
  CLKNV1_8TH40 U170 ( .I(compare_reg[23]), .ZN(n22) );
  CLKNV1_8TH40 U171 ( .I(compare_reg[22]), .ZN(n24) );
  OAI22V0_8TH40 U172 ( .A1(n4), .A2(n26), .B1(n6), .B2(n27), .ZN(n452) );
  OAI22V0_8TH40 U173 ( .A1(n4), .A2(n28), .B1(n6), .B2(n29), .ZN(n451) );
  OAI22V0_8TH40 U174 ( .A1(n4), .A2(n30), .B1(n6), .B2(n31), .ZN(n450) );
  CLKNV1_8TH40 U175 ( .I(compare_reg[18]), .ZN(n32) );
  OAI22V0_8TH40 U176 ( .A1(n4), .A2(n34), .B1(n6), .B2(n35), .ZN(n448) );
  OAI22V0_8TH40 U177 ( .A1(n4), .A2(n36), .B1(n6), .B2(n37), .ZN(n447) );
  OAI22V0_8TH40 U178 ( .A1(n4), .A2(n38), .B1(n6), .B2(n39), .ZN(n446) );
  CLKNV1_8TH40 U179 ( .I(compare_reg[14]), .ZN(n40) );
  CLKNV1_8TH40 U180 ( .I(compare_reg[13]), .ZN(n42) );
  CLKNV1_8TH40 U181 ( .I(compare_reg[12]), .ZN(n44) );
  CLKNV1_8TH40 U182 ( .I(compare_reg[11]), .ZN(n46) );
  CLKNV1_8TH40 U183 ( .I(compare_reg[10]), .ZN(n48) );
  CLKNV1_8TH40 U184 ( .I(compare_reg[9]), .ZN(n50) );
  CLKNV1_8TH40 U185 ( .I(compare_reg[8]), .ZN(n52) );
  OAI22V0_8TH40 U186 ( .A1(n4), .A2(n54), .B1(n6), .B2(n55), .ZN(n438) );
  OAI22V0_8TH40 U187 ( .A1(n4), .A2(n56), .B1(n6), .B2(n57), .ZN(n437) );
  CLKNV1_8TH40 U188 ( .I(compare_reg[5]), .ZN(n58) );
  CLKNV1_8TH40 U189 ( .I(compare_reg[4]), .ZN(n60) );
  CLKNV1_8TH40 U190 ( .I(compare_reg[3]), .ZN(n62) );
  CLKNV1_8TH40 U191 ( .I(compare_reg[2]), .ZN(n64) );
  OAI22V0_8TH40 U192 ( .A1(n4), .A2(n66), .B1(n6), .B2(n67), .ZN(n432) );
  CLKNAND2V1_8TH40 U193 ( .A1(n225), .A2(n4), .ZN(n6) );
  CLKNV1_8TH40 U194 ( .I(compare_reg[0]), .ZN(n68) );
  NOR4V0P5_8TH40 U195 ( .A1(compare_reg[23]), .A2(compare_reg[22]), .A3(
        compare_reg[21]), .A4(compare_reg[20]), .ZN(n77) );
  NOR4V0P5_8TH40 U196 ( .A1(compare_reg[1]), .A2(compare_reg[19]), .A3(
        compare_reg[18]), .A4(compare_reg[17]), .ZN(n76) );
  NOR4V0P5_8TH40 U197 ( .A1(compare_reg[16]), .A2(compare_reg[15]), .A3(
        compare_reg[14]), .A4(compare_reg[13]), .ZN(n75) );
  NOR4V0P5_8TH40 U198 ( .A1(compare_reg[12]), .A2(compare_reg[11]), .A3(
        compare_reg[10]), .A4(compare_reg[0]), .ZN(n74) );
  NOR4V0P5_8TH40 U199 ( .A1(compare_reg[9]), .A2(compare_reg[8]), .A3(
        compare_reg[7]), .A4(compare_reg[6]), .ZN(n81) );
  NOR4V0P5_8TH40 U200 ( .A1(compare_reg[5]), .A2(compare_reg[4]), .A3(
        compare_reg[3]), .A4(compare_reg[31]), .ZN(n80) );
  NOR4V0P5_8TH40 U201 ( .A1(compare_reg[30]), .A2(compare_reg[2]), .A3(
        compare_reg[29]), .A4(compare_reg[28]), .ZN(n79) );
  NOR4V0P5_8TH40 U202 ( .A1(compare_reg[27]), .A2(compare_reg[26]), .A3(
        compare_reg[25]), .A4(compare_reg[24]), .ZN(n78) );
  INAND4V0_8TH40 U203 ( .A1(cp0_reg_waddr[2]), .B1(cp0_reg_waddr[1]), .B2(
        cp0_reg_waddr[0]), .B3(n83), .ZN(n82) );
  OAI22V0_8TH40 U204 ( .A1(n84), .A2(n85), .B1(n7), .B2(n86), .ZN(n429) );
  OAI22V0_8TH40 U205 ( .A1(n84), .A2(n87), .B1(n9), .B2(n86), .ZN(n428) );
  OAI22V0_8TH40 U206 ( .A1(n84), .A2(n88), .B1(n11), .B2(n86), .ZN(n427) );
  NOR2V0P5_8TH40 U207 ( .A1(cp0_reg_wdata[28]), .A2(rst), .ZN(n90) );
  OAI22V0_8TH40 U208 ( .A1(n84), .A2(n91), .B1(n15), .B2(n86), .ZN(n425) );
  OAI22V0_8TH40 U209 ( .A1(n84), .A2(n92), .B1(n17), .B2(n86), .ZN(n424) );
  OAI22V0_8TH40 U210 ( .A1(n84), .A2(n93), .B1(n19), .B2(n86), .ZN(n423) );
  OAI22V0_8TH40 U211 ( .A1(n84), .A2(n94), .B1(n21), .B2(n86), .ZN(n422) );
  OAI22V0_8TH40 U212 ( .A1(n84), .A2(n95), .B1(n23), .B2(n86), .ZN(n421) );
  CLKNV1_8TH40 U213 ( .I(status_reg[22]), .ZN(n96) );
  OAI22V0_8TH40 U214 ( .A1(n84), .A2(n97), .B1(n27), .B2(n86), .ZN(n419) );
  OAI22V0_8TH40 U215 ( .A1(n84), .A2(n98), .B1(n29), .B2(n86), .ZN(n418) );
  OAI22V0_8TH40 U216 ( .A1(n84), .A2(n99), .B1(n31), .B2(n86), .ZN(n417) );
  OAI22V0_8TH40 U217 ( .A1(n84), .A2(n100), .B1(n33), .B2(n86), .ZN(n416) );
  OAI22V0_8TH40 U218 ( .A1(n84), .A2(n101), .B1(n35), .B2(n86), .ZN(n415) );
  OAI22V0_8TH40 U219 ( .A1(n84), .A2(n102), .B1(n37), .B2(n86), .ZN(n414) );
  CLKNV1_8TH40 U220 ( .I(status_reg[15]), .ZN(n103) );
  OAI22V0_8TH40 U221 ( .A1(n84), .A2(n104), .B1(n41), .B2(n86), .ZN(n412) );
  OAI22V0_8TH40 U222 ( .A1(n84), .A2(n105), .B1(n43), .B2(n86), .ZN(n411) );
  OAI22V0_8TH40 U223 ( .A1(n84), .A2(n106), .B1(n45), .B2(n86), .ZN(n410) );
  OAI22V0_8TH40 U224 ( .A1(n84), .A2(n107), .B1(n47), .B2(n86), .ZN(n409) );
  OAI22V0_8TH40 U225 ( .A1(n84), .A2(n108), .B1(n49), .B2(n86), .ZN(n408) );
  OAI22V0_8TH40 U226 ( .A1(n84), .A2(n109), .B1(n51), .B2(n86), .ZN(n407) );
  CLKNV1_8TH40 U227 ( .I(status_reg[8]), .ZN(n110) );
  OAI22V0_8TH40 U228 ( .A1(n84), .A2(n111), .B1(n55), .B2(n86), .ZN(n405) );
  OAI22V0_8TH40 U229 ( .A1(n84), .A2(n112), .B1(n57), .B2(n86), .ZN(n404) );
  OAI22V0_8TH40 U230 ( .A1(n84), .A2(n113), .B1(n59), .B2(n86), .ZN(n403) );
  OAI22V0_8TH40 U231 ( .A1(n84), .A2(n114), .B1(n61), .B2(n86), .ZN(n402) );
  OAI22V0_8TH40 U232 ( .A1(n84), .A2(n115), .B1(n63), .B2(n86), .ZN(n401) );
  OAI22V0_8TH40 U233 ( .A1(n84), .A2(n116), .B1(n65), .B2(n86), .ZN(n400) );
  AOI211V0_8TH40 U234 ( .A1(n120), .A2(n121), .B(n122), .C(n123), .ZN(n119) );
  OAI211V0_8TH40 U235 ( .A1(n125), .A2(n67), .B(n126), .C(n127), .ZN(n124) );
  CLKNV1_8TH40 U236 ( .I(cause_reg[2]), .ZN(n128) );
  CLKNV1_8TH40 U237 ( .I(cause_reg[3]), .ZN(n130) );
  INAND2V0_8TH40 U238 ( .A1(n132), .B1(n120), .ZN(n129) );
  CLKNV1_8TH40 U239 ( .I(cause_reg[4]), .ZN(n133) );
  CLKNAND2V1_8TH40 U240 ( .A1(n122), .A2(n225), .ZN(n132) );
  CLKNV1_8TH40 U241 ( .I(cause_reg[5]), .ZN(n134) );
  NAND3V0P5_8TH40 U242 ( .A1(n126), .A2(n225), .A3(n127), .ZN(n122) );
  MUX2NV0_8TH40 U243 ( .I0(cause_reg[31]), .I1(in_delayslot_i), .S(n136), .ZN(
        n135) );
  AO222V0_8TH40 U244 ( .A1(N290), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[0]), 
        .C1(epc_reg[0]), .C2(n139), .Z(n393) );
  AO222V0_8TH40 U245 ( .A1(N291), .A2(n137), .B1(n138), .B2(cp0_reg_wdata[1]), 
        .C1(epc_reg[1]), .C2(n139), .Z(n392) );
  OA211V0_8TH40 U246 ( .A1(status_reg[1]), .A2(n140), .B(n141), .C(n142), .Z(
        n138) );
  AND2V0_8TH40 U247 ( .A1(n142), .A2(n136), .Z(n137) );
  NOR2V0P5_8TH40 U248 ( .A1(rst), .A2(n139), .ZN(n142) );
  OAI21V0_8TH40 U249 ( .A1(status_reg[1]), .A2(n127), .B(n126), .ZN(n136) );
  NAND4V0P5_8TH40 U250 ( .A1(except_type_i[0]), .A2(n131), .A3(n144), .A4(n145), .ZN(n126) );
  I2NAND4V0_8TH40 U251 ( .A1(n3), .A2(cp0_reg_waddr[0]), .B1(cp0_reg_waddr[1]), 
        .B2(n141), .ZN(n143) );
  INAND2V0_8TH40 U252 ( .A1(n140), .B1(n127), .ZN(n141) );
  AOI32V0_8TH40 U253 ( .A1(except_type_i[3]), .A2(n144), .A3(n121), .B1(n131), 
        .B2(n120), .ZN(n127) );
  CLKNV1_8TH40 U254 ( .I(except_type_i[1]), .ZN(n131) );
  CLKNV1_8TH40 U255 ( .I(except_type_i[0]), .ZN(n121) );
  IOA21V0_8TH40 U256 ( .A1(n120), .A2(except_type_i[1]), .B(n125), .ZN(n140)
         );
  CLKNAND2V1_8TH40 U257 ( .A1(except_type_i[0]), .A2(n144), .ZN(n147) );
  NOR2V0P5_8TH40 U258 ( .A1(n144), .A2(n145), .ZN(n120) );
  CLKNV1_8TH40 U259 ( .I(except_type_i[3]), .ZN(n145) );
  CLKNV1_8TH40 U260 ( .I(except_type_i[2]), .ZN(n144) );
  OAI22V0_8TH40 U261 ( .A1(n84), .A2(n148), .B1(n69), .B2(n86), .ZN(n361) );
  CLKNAND2V1_8TH40 U262 ( .A1(n225), .A2(n84), .ZN(n86) );
  INAND2V0_8TH40 U263 ( .A1(n123), .B1(n225), .ZN(n84) );
  NOR3V0P5_8TH40 U264 ( .A1(cp0_reg_waddr[0]), .A2(cp0_reg_waddr[1]), .A3(n3), 
        .ZN(n123) );
  CLKNAND2V1_8TH40 U265 ( .A1(cp0_reg_waddr[2]), .A2(n83), .ZN(n3) );
  AOI22V0_8TH40 U266 ( .A1(count_reg[31]), .A2(n152), .B1(n153), .B2(
        epc_reg[31]), .ZN(n151) );
  AOI22V0_8TH40 U267 ( .A1(cause_reg[31]), .A2(n154), .B1(n155), .B2(
        compare_reg[31]), .ZN(n150) );
  AOI22V0_8TH40 U268 ( .A1(count_reg[30]), .A2(n152), .B1(n153), .B2(
        epc_reg[30]), .ZN(n157) );
  CLKNV1_8TH40 U269 ( .I(compare_reg[30]), .ZN(n8) );
  AOI22V0_8TH40 U270 ( .A1(count_reg[29]), .A2(n152), .B1(n153), .B2(
        epc_reg[29]), .ZN(n158) );
  CLKNV1_8TH40 U271 ( .I(compare_reg[29]), .ZN(n10) );
  AOI22V0_8TH40 U272 ( .A1(count_reg[28]), .A2(n152), .B1(n153), .B2(
        epc_reg[28]), .ZN(n159) );
  CLKNV1_8TH40 U273 ( .I(compare_reg[28]), .ZN(n12) );
  AOI22V0_8TH40 U274 ( .A1(count_reg[27]), .A2(n152), .B1(n153), .B2(
        epc_reg[27]), .ZN(n160) );
  CLKNV1_8TH40 U275 ( .I(compare_reg[27]), .ZN(n14) );
  AOI22V0_8TH40 U276 ( .A1(count_reg[26]), .A2(n152), .B1(n153), .B2(
        epc_reg[26]), .ZN(n161) );
  CLKNV1_8TH40 U277 ( .I(compare_reg[26]), .ZN(n16) );
  AOI22V0_8TH40 U278 ( .A1(count_reg[25]), .A2(n152), .B1(n153), .B2(
        epc_reg[25]), .ZN(n162) );
  CLKNV1_8TH40 U279 ( .I(compare_reg[25]), .ZN(n18) );
  AOI22V0_8TH40 U280 ( .A1(count_reg[24]), .A2(n152), .B1(n153), .B2(
        epc_reg[24]), .ZN(n164) );
  AOI21V0_8TH40 U281 ( .A1(n155), .A2(compare_reg[24]), .B(n165), .ZN(n163) );
  AOI22V0_8TH40 U282 ( .A1(count_reg[23]), .A2(n152), .B1(n153), .B2(
        epc_reg[23]), .ZN(n167) );
  AOI22V0_8TH40 U283 ( .A1(n172), .A2(status_reg[22]), .B1(count_reg[22]), 
        .B2(n152), .ZN(n170) );
  CLKNV1_8TH40 U284 ( .I(epc_reg[22]), .ZN(n168) );
  AOI22V0_8TH40 U285 ( .A1(count_reg[21]), .A2(n152), .B1(n153), .B2(
        epc_reg[21]), .ZN(n173) );
  CLKNV1_8TH40 U286 ( .I(compare_reg[21]), .ZN(n26) );
  AOI22V0_8TH40 U287 ( .A1(count_reg[20]), .A2(n152), .B1(n153), .B2(
        epc_reg[20]), .ZN(n174) );
  CLKNV1_8TH40 U288 ( .I(compare_reg[20]), .ZN(n28) );
  AOI22V0_8TH40 U289 ( .A1(count_reg[19]), .A2(n152), .B1(n153), .B2(
        epc_reg[19]), .ZN(n175) );
  CLKNV1_8TH40 U290 ( .I(compare_reg[19]), .ZN(n30) );
  AOI22V0_8TH40 U291 ( .A1(count_reg[18]), .A2(n152), .B1(n153), .B2(
        epc_reg[18]), .ZN(n177) );
  AOI21V0_8TH40 U292 ( .A1(n155), .A2(compare_reg[18]), .B(n165), .ZN(n176) );
  AOI22V0_8TH40 U293 ( .A1(count_reg[17]), .A2(n152), .B1(n153), .B2(
        epc_reg[17]), .ZN(n178) );
  CLKNV1_8TH40 U294 ( .I(compare_reg[17]), .ZN(n34) );
  AOI22V0_8TH40 U295 ( .A1(count_reg[16]), .A2(n152), .B1(n153), .B2(
        epc_reg[16]), .ZN(n179) );
  CLKNV1_8TH40 U296 ( .I(compare_reg[16]), .ZN(n36) );
  AOI222V0_8TH40 U297 ( .A1(n153), .A2(epc_reg[15]), .B1(n172), .B2(
        status_reg[15]), .C1(count_reg[15]), .C2(n152), .ZN(n181) );
  CLKNV1_8TH40 U298 ( .I(n184), .ZN(n182) );
  CLKNV1_8TH40 U299 ( .I(compare_reg[15]), .ZN(n38) );
  AOI22V0_8TH40 U300 ( .A1(count_reg[14]), .A2(n152), .B1(n153), .B2(
        epc_reg[14]), .ZN(n186) );
  AOI22V0_8TH40 U301 ( .A1(cause_reg[14]), .A2(n154), .B1(n155), .B2(
        compare_reg[14]), .ZN(n185) );
  CLKNV1_8TH40 U302 ( .I(status_reg[14]), .ZN(n104) );
  AOI22V0_8TH40 U303 ( .A1(count_reg[13]), .A2(n152), .B1(n153), .B2(
        epc_reg[13]), .ZN(n188) );
  AOI22V0_8TH40 U304 ( .A1(cause_reg[13]), .A2(n154), .B1(n155), .B2(
        compare_reg[13]), .ZN(n187) );
  CLKNV1_8TH40 U305 ( .I(status_reg[13]), .ZN(n105) );
  AOI22V0_8TH40 U306 ( .A1(count_reg[12]), .A2(n152), .B1(n153), .B2(
        epc_reg[12]), .ZN(n190) );
  AOI22V0_8TH40 U307 ( .A1(cause_reg[12]), .A2(n154), .B1(n155), .B2(
        compare_reg[12]), .ZN(n189) );
  CLKNV1_8TH40 U308 ( .I(status_reg[12]), .ZN(n106) );
  AOI22V0_8TH40 U309 ( .A1(count_reg[11]), .A2(n152), .B1(n153), .B2(
        epc_reg[11]), .ZN(n192) );
  AOI22V0_8TH40 U310 ( .A1(cause_reg[11]), .A2(n154), .B1(n155), .B2(
        compare_reg[11]), .ZN(n191) );
  CLKNV1_8TH40 U311 ( .I(status_reg[11]), .ZN(n107) );
  AOI22V0_8TH40 U312 ( .A1(count_reg[10]), .A2(n152), .B1(n153), .B2(
        epc_reg[10]), .ZN(n194) );
  AOI22V0_8TH40 U313 ( .A1(cause_reg[10]), .A2(n154), .B1(n155), .B2(
        compare_reg[10]), .ZN(n193) );
  CLKNV1_8TH40 U314 ( .I(status_reg[10]), .ZN(n108) );
  AOI22V0_8TH40 U315 ( .A1(count_reg[9]), .A2(n152), .B1(n153), .B2(epc_reg[9]), .ZN(n196) );
  AOI22V0_8TH40 U316 ( .A1(cause_reg[9]), .A2(n154), .B1(n155), .B2(
        compare_reg[9]), .ZN(n195) );
  CLKNV1_8TH40 U317 ( .I(status_reg[9]), .ZN(n109) );
  AOI221V0_8TH40 U318 ( .A1(n155), .A2(compare_reg[8]), .B1(cause_reg[8]), 
        .B2(n154), .C(n165), .ZN(n199) );
  AOI22V0_8TH40 U319 ( .A1(n172), .A2(status_reg[8]), .B1(count_reg[8]), .B2(
        n152), .ZN(n198) );
  CLKNV1_8TH40 U320 ( .I(n149), .ZN(n172) );
  CLKNV1_8TH40 U321 ( .I(epc_reg[8]), .ZN(n197) );
  AOI22V0_8TH40 U322 ( .A1(count_reg[7]), .A2(n152), .B1(n153), .B2(epc_reg[7]), .ZN(n200) );
  CLKNV1_8TH40 U323 ( .I(compare_reg[7]), .ZN(n54) );
  AOI22V0_8TH40 U324 ( .A1(count_reg[6]), .A2(n152), .B1(n153), .B2(epc_reg[6]), .ZN(n201) );
  CLKNV1_8TH40 U325 ( .I(compare_reg[6]), .ZN(n56) );
  AOI22V0_8TH40 U326 ( .A1(count_reg[5]), .A2(n152), .B1(n153), .B2(epc_reg[5]), .ZN(n203) );
  AOI22V0_8TH40 U327 ( .A1(n154), .A2(cause_reg[5]), .B1(n155), .B2(
        compare_reg[5]), .ZN(n202) );
  AOI22V0_8TH40 U328 ( .A1(count_reg[4]), .A2(n152), .B1(n153), .B2(epc_reg[4]), .ZN(n205) );
  AOI22V0_8TH40 U329 ( .A1(n154), .A2(cause_reg[4]), .B1(n155), .B2(
        compare_reg[4]), .ZN(n204) );
  AOI22V0_8TH40 U330 ( .A1(count_reg[3]), .A2(n152), .B1(n153), .B2(epc_reg[3]), .ZN(n207) );
  AOI22V0_8TH40 U331 ( .A1(n154), .A2(cause_reg[3]), .B1(n155), .B2(
        compare_reg[3]), .ZN(n206) );
  AOI22V0_8TH40 U332 ( .A1(count_reg[2]), .A2(n152), .B1(n153), .B2(epc_reg[2]), .ZN(n209) );
  AOI22V0_8TH40 U333 ( .A1(n154), .A2(cause_reg[2]), .B1(n155), .B2(
        compare_reg[2]), .ZN(n208) );
  I2NOR3V1_8TH40 U334 ( .A1(n210), .A2(n183), .B(n211), .ZN(n154) );
  AOI22V0_8TH40 U335 ( .A1(count_reg[1]), .A2(n152), .B1(n153), .B2(epc_reg[1]), .ZN(n212) );
  CLKNV1_8TH40 U336 ( .I(status_reg[1]), .ZN(n118) );
  CLKNV1_8TH40 U337 ( .I(compare_reg[1]), .ZN(n66) );
  AOI22V0_8TH40 U338 ( .A1(count_reg[0]), .A2(n152), .B1(n153), .B2(epc_reg[0]), .ZN(n214) );
  CLKNV1_8TH40 U339 ( .I(n169), .ZN(n153) );
  CLKNAND2V1_8TH40 U340 ( .A1(n215), .A2(n216), .ZN(n169) );
  I2NOR3V1_8TH40 U341 ( .A1(n183), .A2(n210), .B(cp0_reg_raddr[2]), .ZN(n152)
         );
  AOI21V0_8TH40 U342 ( .A1(n155), .A2(compare_reg[0]), .B(n165), .ZN(n213) );
  I2NOR3V1_8TH40 U343 ( .A1(n216), .A2(n210), .B(n211), .ZN(n165) );
  CLKNV1_8TH40 U344 ( .I(n156), .ZN(n155) );
  NAND3V0P5_8TH40 U345 ( .A1(n210), .A2(n211), .A3(n216), .ZN(n156) );
  INOR2V0_8TH40 U346 ( .A1(cp0_reg_raddr[1]), .B1(rst), .ZN(n216) );
  CLKNAND2V1_8TH40 U347 ( .A1(n215), .A2(n183), .ZN(n149) );
  NOR2V0P5_8TH40 U348 ( .A1(cp0_reg_raddr[1]), .A2(rst), .ZN(n183) );
  CLKNV1_8TH40 U349 ( .I(status_reg[0]), .ZN(n148) );
  OAI211V0_8TH40 U350 ( .A1(cp0_reg_raddr[1]), .A2(n184), .B(n217), .C(n218), 
        .ZN(N867) );
  NOR2V0P5_8TH40 U351 ( .A1(rst), .A2(n210), .ZN(n218) );
  NOR3V0P5_8TH40 U352 ( .A1(n219), .A2(cp0_reg_raddr[4]), .A3(n220), .ZN(n210)
         );
  CLKNV1_8TH40 U353 ( .I(n215), .ZN(n217) );
  NOR4V0P5_8TH40 U354 ( .A1(n211), .A2(n220), .A3(cp0_reg_raddr[0]), .A4(
        cp0_reg_raddr[4]), .ZN(n215) );
  NAND4V0P5_8TH40 U355 ( .A1(cp0_reg_raddr[4]), .A2(n219), .A3(n211), .A4(n220), .ZN(n184) );
  CLKNV1_8TH40 U356 ( .I(cp0_reg_raddr[2]), .ZN(n211) );
  CLKNV1_8TH40 U357 ( .I(cp0_reg_raddr[0]), .ZN(n219) );
  CLKNV1_8TH40 U358 ( .I(cp0_reg_wdata[31]), .ZN(n7) );
  CLKNV1_8TH40 U359 ( .I(cp0_reg_wdata[30]), .ZN(n9) );
  CLKNV1_8TH40 U360 ( .I(cp0_reg_wdata[29]), .ZN(n11) );
  CLKNV1_8TH40 U361 ( .I(cp0_reg_wdata[28]), .ZN(n13) );
  CLKNV1_8TH40 U362 ( .I(cp0_reg_wdata[27]), .ZN(n15) );
  CLKNV1_8TH40 U363 ( .I(cp0_reg_wdata[26]), .ZN(n17) );
  CLKNV1_8TH40 U364 ( .I(cp0_reg_wdata[25]), .ZN(n19) );
  CLKNV1_8TH40 U365 ( .I(cp0_reg_wdata[24]), .ZN(n21) );
  CLKNV1_8TH40 U366 ( .I(cp0_reg_wdata[23]), .ZN(n23) );
  CLKNV1_8TH40 U367 ( .I(cp0_reg_wdata[22]), .ZN(n25) );
  CLKNV1_8TH40 U368 ( .I(cp0_reg_wdata[21]), .ZN(n27) );
  CLKNV1_8TH40 U369 ( .I(cp0_reg_wdata[20]), .ZN(n29) );
  CLKNV1_8TH40 U370 ( .I(cp0_reg_wdata[19]), .ZN(n31) );
  CLKNV1_8TH40 U371 ( .I(cp0_reg_wdata[18]), .ZN(n33) );
  CLKNV1_8TH40 U372 ( .I(cp0_reg_wdata[17]), .ZN(n35) );
  CLKNV1_8TH40 U373 ( .I(cp0_reg_wdata[16]), .ZN(n37) );
  CLKNV1_8TH40 U374 ( .I(cp0_reg_wdata[15]), .ZN(n39) );
  CLKNV1_8TH40 U375 ( .I(cp0_reg_wdata[14]), .ZN(n41) );
  CLKNV1_8TH40 U376 ( .I(cp0_reg_wdata[13]), .ZN(n43) );
  CLKNV1_8TH40 U377 ( .I(cp0_reg_wdata[12]), .ZN(n45) );
  CLKNV1_8TH40 U378 ( .I(cp0_reg_wdata[11]), .ZN(n47) );
  CLKNV1_8TH40 U379 ( .I(cp0_reg_wdata[10]), .ZN(n49) );
  CLKNV1_8TH40 U380 ( .I(cp0_reg_wdata[9]), .ZN(n51) );
  CLKNV1_8TH40 U381 ( .I(cp0_reg_wdata[8]), .ZN(n53) );
  CLKNV1_8TH40 U382 ( .I(cp0_reg_wdata[7]), .ZN(n55) );
  CLKNV1_8TH40 U383 ( .I(cp0_reg_wdata[6]), .ZN(n57) );
  CLKNV1_8TH40 U384 ( .I(cp0_reg_wdata[5]), .ZN(n59) );
  CLKNV1_8TH40 U385 ( .I(cp0_reg_wdata[4]), .ZN(n61) );
  CLKNV1_8TH40 U386 ( .I(cp0_reg_wdata[3]), .ZN(n63) );
  CLKNV1_8TH40 U387 ( .I(cp0_reg_wdata[2]), .ZN(n65) );
  CLKNV1_8TH40 U388 ( .I(cp0_reg_wdata[1]), .ZN(n67) );
  NOR2V0P5_8TH40 U389 ( .A1(n223), .A2(rst), .ZN(n222) );
  CLKNAND2V1_8TH40 U390 ( .A1(n223), .A2(n225), .ZN(n221) );
  CLKNV1_8TH40 U391 ( .I(rst), .ZN(n225) );
  I2NOR4V0_8TH40 U392 ( .A1(n83), .A2(cp0_reg_waddr[0]), .B1(cp0_reg_waddr[1]), 
        .B2(cp0_reg_waddr[2]), .ZN(n223) );
  I2NOR3V1_8TH40 U393 ( .A1(cp0_reg_we), .A2(cp0_reg_waddr[3]), .B(
        cp0_reg_waddr[4]), .ZN(n83) );
  CLKNV1_8TH40 U394 ( .I(cp0_reg_wdata[0]), .ZN(n69) );
endmodule


module wb_interface_0 ( clk, rst, stall_ctrl, cpu_ce_i, cpu_data_i, cpu_addr_i, 
        cpu_we_i, cpu_sel_i, cpu_data_o, wb_data_i, wb_ack_i, wb_addr_o, 
        wb_data_o, wb_we_o, wb_sel_o, wb_stb_o, wb_cyc_o, stall_req, 
        flush_i_BAR );
  input [5:0] stall_ctrl;
  input [31:0] cpu_data_i;
  input [31:0] cpu_addr_i;
  input [3:0] cpu_sel_i;
  output [31:0] cpu_data_o;
  input [31:0] wb_data_i;
  output [31:0] wb_addr_o;
  output [31:0] wb_data_o;
  output [3:0] wb_sel_o;
  input clk, rst, cpu_ce_i, cpu_we_i, wb_ack_i, flush_i_BAR;
  output wb_we_o, wb_stb_o, wb_cyc_o, stall_req;
  wire   N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n1, n2, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86;
  wire   [1:0] wb_state;

  DQV4_8TH40 wb_state_reg_0_ ( .D(n195), .CK(clk), .Q(wb_state[0]) );
  DQV4_8TH40 wb_state_reg_1_ ( .D(n194), .CK(clk), .Q(wb_state[1]) );
  DQNV4_8TH40 data_buf_reg_31_ ( .D(n162), .CK(clk), .QN(n3) );
  DQNV4_8TH40 data_buf_reg_30_ ( .D(n163), .CK(clk), .QN(n4) );
  DQNV4_8TH40 data_buf_reg_29_ ( .D(n164), .CK(clk), .QN(n5) );
  DQNV4_8TH40 data_buf_reg_28_ ( .D(n165), .CK(clk), .QN(n6) );
  DQNV4_8TH40 data_buf_reg_27_ ( .D(n166), .CK(clk), .QN(n7) );
  DQNV4_8TH40 data_buf_reg_26_ ( .D(n167), .CK(clk), .QN(n8) );
  DQNV4_8TH40 data_buf_reg_25_ ( .D(n168), .CK(clk), .QN(n9) );
  DQNV4_8TH40 data_buf_reg_24_ ( .D(n169), .CK(clk), .QN(n10) );
  DQNV4_8TH40 data_buf_reg_23_ ( .D(n170), .CK(clk), .QN(n11) );
  DQNV4_8TH40 data_buf_reg_22_ ( .D(n171), .CK(clk), .QN(n12) );
  DQNV4_8TH40 data_buf_reg_21_ ( .D(n172), .CK(clk), .QN(n13) );
  DQNV4_8TH40 data_buf_reg_20_ ( .D(n173), .CK(clk), .QN(n14) );
  DQNV4_8TH40 data_buf_reg_19_ ( .D(n174), .CK(clk), .QN(n15) );
  DQNV4_8TH40 data_buf_reg_18_ ( .D(n175), .CK(clk), .QN(n16) );
  DQNV4_8TH40 data_buf_reg_17_ ( .D(n176), .CK(clk), .QN(n17) );
  DQNV4_8TH40 data_buf_reg_16_ ( .D(n177), .CK(clk), .QN(n18) );
  DQNV4_8TH40 data_buf_reg_15_ ( .D(n178), .CK(clk), .QN(n19) );
  DQNV4_8TH40 data_buf_reg_14_ ( .D(n179), .CK(clk), .QN(n20) );
  DQNV4_8TH40 data_buf_reg_13_ ( .D(n180), .CK(clk), .QN(n21) );
  DQNV4_8TH40 data_buf_reg_12_ ( .D(n181), .CK(clk), .QN(n22) );
  DQNV4_8TH40 data_buf_reg_11_ ( .D(n182), .CK(clk), .QN(n23) );
  DQNV4_8TH40 data_buf_reg_10_ ( .D(n183), .CK(clk), .QN(n24) );
  DQNV4_8TH40 data_buf_reg_9_ ( .D(n184), .CK(clk), .QN(n25) );
  DQNV4_8TH40 data_buf_reg_8_ ( .D(n185), .CK(clk), .QN(n26) );
  DQNV4_8TH40 data_buf_reg_7_ ( .D(n186), .CK(clk), .QN(n27) );
  DQNV4_8TH40 data_buf_reg_6_ ( .D(n187), .CK(clk), .QN(n28) );
  DQNV4_8TH40 data_buf_reg_5_ ( .D(n188), .CK(clk), .QN(n29) );
  DQNV4_8TH40 data_buf_reg_4_ ( .D(n189), .CK(clk), .QN(n30) );
  DQNV4_8TH40 data_buf_reg_3_ ( .D(n190), .CK(clk), .QN(n31) );
  DQNV4_8TH40 data_buf_reg_2_ ( .D(n191), .CK(clk), .QN(n32) );
  DQNV4_8TH40 data_buf_reg_1_ ( .D(n192), .CK(clk), .QN(n33) );
  DQNV4_8TH40 data_buf_reg_0_ ( .D(n193), .CK(clk), .QN(n34) );
  DQV4_8TH40 wb_sel_o_reg_3_ ( .D(n125), .CK(clk), .Q(wb_sel_o[3]) );
  DQV4_8TH40 wb_sel_o_reg_2_ ( .D(n126), .CK(clk), .Q(wb_sel_o[2]) );
  DQV4_8TH40 wb_sel_o_reg_1_ ( .D(n127), .CK(clk), .Q(wb_sel_o[1]) );
  DQV4_8TH40 wb_sel_o_reg_0_ ( .D(n128), .CK(clk), .Q(wb_sel_o[0]) );
  DQV4_8TH40 wb_we_o_reg ( .D(n129), .CK(clk), .Q(wb_we_o) );
  DQV4_8TH40 wb_data_o_reg_31_ ( .D(n130), .CK(clk), .Q(wb_data_o[31]) );
  DQV4_8TH40 wb_data_o_reg_30_ ( .D(n131), .CK(clk), .Q(wb_data_o[30]) );
  DQV4_8TH40 wb_data_o_reg_29_ ( .D(n132), .CK(clk), .Q(wb_data_o[29]) );
  DQV4_8TH40 wb_data_o_reg_28_ ( .D(n133), .CK(clk), .Q(wb_data_o[28]) );
  DQV4_8TH40 wb_data_o_reg_27_ ( .D(n134), .CK(clk), .Q(wb_data_o[27]) );
  DQV4_8TH40 wb_data_o_reg_26_ ( .D(n135), .CK(clk), .Q(wb_data_o[26]) );
  DQV4_8TH40 wb_data_o_reg_25_ ( .D(n136), .CK(clk), .Q(wb_data_o[25]) );
  DQV4_8TH40 wb_data_o_reg_24_ ( .D(n137), .CK(clk), .Q(wb_data_o[24]) );
  DQV4_8TH40 wb_data_o_reg_23_ ( .D(n138), .CK(clk), .Q(wb_data_o[23]) );
  DQV4_8TH40 wb_data_o_reg_22_ ( .D(n139), .CK(clk), .Q(wb_data_o[22]) );
  DQV4_8TH40 wb_data_o_reg_21_ ( .D(n140), .CK(clk), .Q(wb_data_o[21]) );
  DQV4_8TH40 wb_data_o_reg_20_ ( .D(n141), .CK(clk), .Q(wb_data_o[20]) );
  DQV4_8TH40 wb_data_o_reg_19_ ( .D(n142), .CK(clk), .Q(wb_data_o[19]) );
  DQV4_8TH40 wb_data_o_reg_18_ ( .D(n143), .CK(clk), .Q(wb_data_o[18]) );
  DQV4_8TH40 wb_data_o_reg_17_ ( .D(n144), .CK(clk), .Q(wb_data_o[17]) );
  DQV4_8TH40 wb_data_o_reg_16_ ( .D(n145), .CK(clk), .Q(wb_data_o[16]) );
  DQV4_8TH40 wb_data_o_reg_15_ ( .D(n146), .CK(clk), .Q(wb_data_o[15]) );
  DQV4_8TH40 wb_data_o_reg_14_ ( .D(n147), .CK(clk), .Q(wb_data_o[14]) );
  DQV4_8TH40 wb_data_o_reg_13_ ( .D(n148), .CK(clk), .Q(wb_data_o[13]) );
  DQV4_8TH40 wb_data_o_reg_12_ ( .D(n149), .CK(clk), .Q(wb_data_o[12]) );
  DQV4_8TH40 wb_data_o_reg_11_ ( .D(n150), .CK(clk), .Q(wb_data_o[11]) );
  DQV4_8TH40 wb_data_o_reg_10_ ( .D(n151), .CK(clk), .Q(wb_data_o[10]) );
  DQV4_8TH40 wb_data_o_reg_9_ ( .D(n152), .CK(clk), .Q(wb_data_o[9]) );
  DQV4_8TH40 wb_data_o_reg_8_ ( .D(n153), .CK(clk), .Q(wb_data_o[8]) );
  DQV4_8TH40 wb_data_o_reg_7_ ( .D(n154), .CK(clk), .Q(wb_data_o[7]) );
  DQV4_8TH40 wb_data_o_reg_6_ ( .D(n155), .CK(clk), .Q(wb_data_o[6]) );
  DQV4_8TH40 wb_data_o_reg_5_ ( .D(n156), .CK(clk), .Q(wb_data_o[5]) );
  DQV4_8TH40 wb_data_o_reg_4_ ( .D(n157), .CK(clk), .Q(wb_data_o[4]) );
  DQV4_8TH40 wb_data_o_reg_3_ ( .D(n158), .CK(clk), .Q(wb_data_o[3]) );
  DQV4_8TH40 wb_data_o_reg_2_ ( .D(n159), .CK(clk), .Q(wb_data_o[2]) );
  DQV4_8TH40 wb_data_o_reg_1_ ( .D(n160), .CK(clk), .Q(wb_data_o[1]) );
  DQV4_8TH40 wb_data_o_reg_0_ ( .D(n161), .CK(clk), .Q(wb_data_o[0]) );
  DQV4_8TH40 wb_addr_o_reg_31_ ( .D(n124), .CK(clk), .Q(wb_addr_o[31]) );
  DQV4_8TH40 wb_addr_o_reg_30_ ( .D(n123), .CK(clk), .Q(wb_addr_o[30]) );
  DQV4_8TH40 wb_addr_o_reg_29_ ( .D(n122), .CK(clk), .Q(wb_addr_o[29]) );
  DQV4_8TH40 wb_addr_o_reg_28_ ( .D(n121), .CK(clk), .Q(wb_addr_o[28]) );
  DQV4_8TH40 wb_addr_o_reg_27_ ( .D(n120), .CK(clk), .Q(wb_addr_o[27]) );
  DQV4_8TH40 wb_addr_o_reg_26_ ( .D(n119), .CK(clk), .Q(wb_addr_o[26]) );
  DQV4_8TH40 wb_addr_o_reg_25_ ( .D(n118), .CK(clk), .Q(wb_addr_o[25]) );
  DQV4_8TH40 wb_addr_o_reg_24_ ( .D(n117), .CK(clk), .Q(wb_addr_o[24]) );
  DQV4_8TH40 wb_addr_o_reg_23_ ( .D(n116), .CK(clk), .Q(wb_addr_o[23]) );
  DQV4_8TH40 wb_addr_o_reg_22_ ( .D(n115), .CK(clk), .Q(wb_addr_o[22]) );
  DQV4_8TH40 wb_addr_o_reg_21_ ( .D(n114), .CK(clk), .Q(wb_addr_o[21]) );
  DQV4_8TH40 wb_addr_o_reg_20_ ( .D(n113), .CK(clk), .Q(wb_addr_o[20]) );
  DQV4_8TH40 wb_addr_o_reg_19_ ( .D(n112), .CK(clk), .Q(wb_addr_o[19]) );
  DQV4_8TH40 wb_addr_o_reg_18_ ( .D(n111), .CK(clk), .Q(wb_addr_o[18]) );
  DQV4_8TH40 wb_addr_o_reg_17_ ( .D(n110), .CK(clk), .Q(wb_addr_o[17]) );
  DQV4_8TH40 wb_addr_o_reg_16_ ( .D(n109), .CK(clk), .Q(wb_addr_o[16]) );
  DQV4_8TH40 wb_addr_o_reg_15_ ( .D(n108), .CK(clk), .Q(wb_addr_o[15]) );
  DQV4_8TH40 wb_addr_o_reg_14_ ( .D(n107), .CK(clk), .Q(wb_addr_o[14]) );
  DQV4_8TH40 wb_addr_o_reg_13_ ( .D(n106), .CK(clk), .Q(wb_addr_o[13]) );
  DQV4_8TH40 wb_addr_o_reg_12_ ( .D(n105), .CK(clk), .Q(wb_addr_o[12]) );
  DQV4_8TH40 wb_addr_o_reg_11_ ( .D(n104), .CK(clk), .Q(wb_addr_o[11]) );
  DQV4_8TH40 wb_addr_o_reg_10_ ( .D(n103), .CK(clk), .Q(wb_addr_o[10]) );
  DQV4_8TH40 wb_addr_o_reg_9_ ( .D(n102), .CK(clk), .Q(wb_addr_o[9]) );
  DQV4_8TH40 wb_addr_o_reg_8_ ( .D(n101), .CK(clk), .Q(wb_addr_o[8]) );
  DQV4_8TH40 wb_addr_o_reg_7_ ( .D(n100), .CK(clk), .Q(wb_addr_o[7]) );
  DQV4_8TH40 wb_addr_o_reg_6_ ( .D(n99), .CK(clk), .Q(wb_addr_o[6]) );
  DQV4_8TH40 wb_addr_o_reg_5_ ( .D(n98), .CK(clk), .Q(wb_addr_o[5]) );
  DQV4_8TH40 wb_addr_o_reg_4_ ( .D(n97), .CK(clk), .Q(wb_addr_o[4]) );
  DQV4_8TH40 wb_addr_o_reg_3_ ( .D(n96), .CK(clk), .Q(wb_addr_o[3]) );
  DQV4_8TH40 wb_addr_o_reg_2_ ( .D(n95), .CK(clk), .Q(wb_addr_o[2]) );
  DQV4_8TH40 wb_addr_o_reg_1_ ( .D(n94), .CK(clk), .Q(wb_addr_o[1]) );
  DQV4_8TH40 wb_addr_o_reg_0_ ( .D(n93), .CK(clk), .Q(wb_addr_o[0]) );
  LAHQV1_8TH40 cpu_data_o_reg_31_ ( .E(N387), .D(N419), .Q(cpu_data_o[31]) );
  LAHQV1_8TH40 cpu_data_o_reg_30_ ( .E(N387), .D(N418), .Q(cpu_data_o[30]) );
  LAHQV1_8TH40 cpu_data_o_reg_29_ ( .E(N387), .D(N417), .Q(cpu_data_o[29]) );
  LAHQV1_8TH40 cpu_data_o_reg_28_ ( .E(N387), .D(N416), .Q(cpu_data_o[28]) );
  LAHQV1_8TH40 cpu_data_o_reg_27_ ( .E(N387), .D(N415), .Q(cpu_data_o[27]) );
  LAHQV1_8TH40 cpu_data_o_reg_26_ ( .E(N387), .D(N414), .Q(cpu_data_o[26]) );
  LAHQV1_8TH40 cpu_data_o_reg_25_ ( .E(N387), .D(N413), .Q(cpu_data_o[25]) );
  LAHQV1_8TH40 cpu_data_o_reg_24_ ( .E(N387), .D(N412), .Q(cpu_data_o[24]) );
  LAHQV1_8TH40 cpu_data_o_reg_23_ ( .E(N387), .D(N411), .Q(cpu_data_o[23]) );
  LAHQV1_8TH40 cpu_data_o_reg_22_ ( .E(N387), .D(N410), .Q(cpu_data_o[22]) );
  LAHQV1_8TH40 cpu_data_o_reg_21_ ( .E(N387), .D(N409), .Q(cpu_data_o[21]) );
  LAHQV1_8TH40 cpu_data_o_reg_20_ ( .E(N387), .D(N408), .Q(cpu_data_o[20]) );
  LAHQV1_8TH40 cpu_data_o_reg_19_ ( .E(N387), .D(N407), .Q(cpu_data_o[19]) );
  LAHQV1_8TH40 cpu_data_o_reg_18_ ( .E(N387), .D(N406), .Q(cpu_data_o[18]) );
  LAHQV1_8TH40 cpu_data_o_reg_17_ ( .E(N387), .D(N405), .Q(cpu_data_o[17]) );
  LAHQV1_8TH40 cpu_data_o_reg_16_ ( .E(N387), .D(N404), .Q(cpu_data_o[16]) );
  LAHQV1_8TH40 cpu_data_o_reg_15_ ( .E(N387), .D(N403), .Q(cpu_data_o[15]) );
  LAHQV1_8TH40 cpu_data_o_reg_14_ ( .E(N387), .D(N402), .Q(cpu_data_o[14]) );
  LAHQV1_8TH40 cpu_data_o_reg_13_ ( .E(N387), .D(N401), .Q(cpu_data_o[13]) );
  LAHQV1_8TH40 cpu_data_o_reg_12_ ( .E(N387), .D(N400), .Q(cpu_data_o[12]) );
  LAHQV1_8TH40 cpu_data_o_reg_11_ ( .E(N387), .D(N399), .Q(cpu_data_o[11]) );
  LAHQV1_8TH40 cpu_data_o_reg_10_ ( .E(N387), .D(N398), .Q(cpu_data_o[10]) );
  LAHQV1_8TH40 cpu_data_o_reg_9_ ( .E(N387), .D(N397), .Q(cpu_data_o[9]) );
  LAHQV1_8TH40 cpu_data_o_reg_8_ ( .E(N387), .D(N396), .Q(cpu_data_o[8]) );
  LAHQV1_8TH40 cpu_data_o_reg_7_ ( .E(N387), .D(N395), .Q(cpu_data_o[7]) );
  LAHQV1_8TH40 cpu_data_o_reg_6_ ( .E(N387), .D(N394), .Q(cpu_data_o[6]) );
  LAHQV1_8TH40 cpu_data_o_reg_5_ ( .E(N387), .D(N393), .Q(cpu_data_o[5]) );
  LAHQV1_8TH40 cpu_data_o_reg_4_ ( .E(N387), .D(N392), .Q(cpu_data_o[4]) );
  LAHQV1_8TH40 cpu_data_o_reg_3_ ( .E(N387), .D(N391), .Q(cpu_data_o[3]) );
  LAHQV1_8TH40 cpu_data_o_reg_2_ ( .E(N387), .D(N390), .Q(cpu_data_o[2]) );
  LAHQV1_8TH40 cpu_data_o_reg_1_ ( .E(N387), .D(N389), .Q(cpu_data_o[1]) );
  LAHQV1_8TH40 cpu_data_o_reg_0_ ( .E(N387), .D(N388), .Q(cpu_data_o[0]) );
  EDQV2_8TH40 wb_cyc_o_reg ( .D(n86), .E(n85), .CK(clk), .Q(wb_cyc_o) );
  EDQV2_8TH40 wb_stb_o_reg ( .D(n86), .E(n85), .CK(clk), .Q(wb_stb_o) );
  AO22V4_8TH40 U3 ( .A1(wb_addr_o[6]), .A2(n36), .B1(cpu_addr_i[6]), .B2(n37), 
        .Z(n99) );
  AO22V4_8TH40 U4 ( .A1(wb_addr_o[5]), .A2(n36), .B1(cpu_addr_i[5]), .B2(n37), 
        .Z(n98) );
  AO22V4_8TH40 U5 ( .A1(wb_addr_o[4]), .A2(n36), .B1(cpu_addr_i[4]), .B2(n37), 
        .Z(n97) );
  AO22V4_8TH40 U6 ( .A1(wb_addr_o[3]), .A2(n36), .B1(cpu_addr_i[3]), .B2(n37), 
        .Z(n96) );
  AO22V4_8TH40 U7 ( .A1(wb_addr_o[2]), .A2(n36), .B1(cpu_addr_i[2]), .B2(n37), 
        .Z(n95) );
  AO22V4_8TH40 U8 ( .A1(wb_addr_o[1]), .A2(n36), .B1(cpu_addr_i[1]), .B2(n37), 
        .Z(n94) );
  AO22V4_8TH40 U9 ( .A1(wb_addr_o[0]), .A2(n36), .B1(cpu_addr_i[0]), .B2(n37), 
        .Z(n93) );
  AO22V4_8TH40 U10 ( .A1(wb_data_o[0]), .A2(n36), .B1(cpu_data_i[0]), .B2(n37), 
        .Z(n161) );
  AO22V4_8TH40 U11 ( .A1(wb_data_o[1]), .A2(n36), .B1(cpu_data_i[1]), .B2(n37), 
        .Z(n160) );
  AO22V4_8TH40 U12 ( .A1(wb_data_o[2]), .A2(n36), .B1(cpu_data_i[2]), .B2(n37), 
        .Z(n159) );
  AO22V4_8TH40 U13 ( .A1(wb_data_o[3]), .A2(n36), .B1(cpu_data_i[3]), .B2(n37), 
        .Z(n158) );
  AO22V4_8TH40 U14 ( .A1(wb_data_o[4]), .A2(n36), .B1(cpu_data_i[4]), .B2(n37), 
        .Z(n157) );
  AO22V4_8TH40 U15 ( .A1(wb_data_o[5]), .A2(n36), .B1(cpu_data_i[5]), .B2(n37), 
        .Z(n156) );
  AO22V4_8TH40 U16 ( .A1(wb_data_o[6]), .A2(n36), .B1(cpu_data_i[6]), .B2(n37), 
        .Z(n155) );
  AO22V4_8TH40 U17 ( .A1(wb_data_o[7]), .A2(n36), .B1(cpu_data_i[7]), .B2(n37), 
        .Z(n154) );
  AO22V4_8TH40 U18 ( .A1(wb_data_o[8]), .A2(n36), .B1(cpu_data_i[8]), .B2(n37), 
        .Z(n153) );
  AO22V4_8TH40 U19 ( .A1(wb_data_o[9]), .A2(n36), .B1(cpu_data_i[9]), .B2(n37), 
        .Z(n152) );
  AO22V4_8TH40 U20 ( .A1(wb_data_o[10]), .A2(n36), .B1(cpu_data_i[10]), .B2(
        n37), .Z(n151) );
  AO22V4_8TH40 U21 ( .A1(wb_data_o[11]), .A2(n36), .B1(cpu_data_i[11]), .B2(
        n37), .Z(n150) );
  AO22V4_8TH40 U22 ( .A1(wb_data_o[12]), .A2(n36), .B1(cpu_data_i[12]), .B2(
        n37), .Z(n149) );
  AO22V4_8TH40 U23 ( .A1(wb_data_o[13]), .A2(n36), .B1(cpu_data_i[13]), .B2(
        n37), .Z(n148) );
  AO22V4_8TH40 U24 ( .A1(wb_data_o[14]), .A2(n36), .B1(cpu_data_i[14]), .B2(
        n37), .Z(n147) );
  AO22V4_8TH40 U25 ( .A1(wb_data_o[15]), .A2(n36), .B1(cpu_data_i[15]), .B2(
        n37), .Z(n146) );
  AO22V4_8TH40 U26 ( .A1(wb_data_o[16]), .A2(n36), .B1(cpu_data_i[16]), .B2(
        n37), .Z(n145) );
  AO22V4_8TH40 U27 ( .A1(wb_data_o[17]), .A2(n36), .B1(cpu_data_i[17]), .B2(
        n37), .Z(n144) );
  AO22V4_8TH40 U28 ( .A1(wb_data_o[18]), .A2(n36), .B1(cpu_data_i[18]), .B2(
        n37), .Z(n143) );
  AO22V4_8TH40 U29 ( .A1(wb_data_o[19]), .A2(n36), .B1(cpu_data_i[19]), .B2(
        n37), .Z(n142) );
  AO22V4_8TH40 U30 ( .A1(wb_data_o[20]), .A2(n36), .B1(cpu_data_i[20]), .B2(
        n37), .Z(n141) );
  AO22V4_8TH40 U31 ( .A1(wb_data_o[21]), .A2(n36), .B1(cpu_data_i[21]), .B2(
        n37), .Z(n140) );
  AO22V4_8TH40 U32 ( .A1(wb_data_o[22]), .A2(n36), .B1(cpu_data_i[22]), .B2(
        n37), .Z(n139) );
  AO22V4_8TH40 U33 ( .A1(wb_data_o[23]), .A2(n36), .B1(cpu_data_i[23]), .B2(
        n37), .Z(n138) );
  AO22V4_8TH40 U34 ( .A1(wb_data_o[24]), .A2(n36), .B1(cpu_data_i[24]), .B2(
        n37), .Z(n137) );
  AO22V4_8TH40 U35 ( .A1(wb_data_o[25]), .A2(n36), .B1(cpu_data_i[25]), .B2(
        n37), .Z(n136) );
  AO22V4_8TH40 U36 ( .A1(wb_data_o[26]), .A2(n36), .B1(cpu_data_i[26]), .B2(
        n37), .Z(n135) );
  AO22V4_8TH40 U37 ( .A1(wb_data_o[27]), .A2(n36), .B1(cpu_data_i[27]), .B2(
        n37), .Z(n134) );
  AO22V4_8TH40 U38 ( .A1(wb_data_o[28]), .A2(n36), .B1(cpu_data_i[28]), .B2(
        n37), .Z(n133) );
  AO22V4_8TH40 U39 ( .A1(wb_data_o[29]), .A2(n36), .B1(cpu_data_i[29]), .B2(
        n37), .Z(n132) );
  AO22V4_8TH40 U40 ( .A1(wb_data_o[30]), .A2(n36), .B1(cpu_data_i[30]), .B2(
        n37), .Z(n131) );
  AO22V4_8TH40 U41 ( .A1(wb_data_o[31]), .A2(n36), .B1(cpu_data_i[31]), .B2(
        n37), .Z(n130) );
  AO22V4_8TH40 U42 ( .A1(wb_sel_o[0]), .A2(n36), .B1(cpu_sel_i[0]), .B2(n37), 
        .Z(n128) );
  AO22V4_8TH40 U43 ( .A1(wb_sel_o[1]), .A2(n36), .B1(cpu_sel_i[1]), .B2(n37), 
        .Z(n127) );
  AO22V4_8TH40 U44 ( .A1(wb_sel_o[2]), .A2(n36), .B1(cpu_sel_i[2]), .B2(n37), 
        .Z(n126) );
  AO22V4_8TH40 U45 ( .A1(wb_sel_o[3]), .A2(n36), .B1(cpu_sel_i[3]), .B2(n37), 
        .Z(n125) );
  AO22V4_8TH40 U46 ( .A1(wb_addr_o[31]), .A2(n36), .B1(cpu_addr_i[31]), .B2(
        n37), .Z(n124) );
  AO22V4_8TH40 U47 ( .A1(wb_addr_o[30]), .A2(n36), .B1(cpu_addr_i[30]), .B2(
        n37), .Z(n123) );
  AO22V4_8TH40 U48 ( .A1(wb_addr_o[29]), .A2(n36), .B1(cpu_addr_i[29]), .B2(
        n37), .Z(n122) );
  AO22V4_8TH40 U49 ( .A1(wb_addr_o[28]), .A2(n36), .B1(cpu_addr_i[28]), .B2(
        n37), .Z(n121) );
  AO22V4_8TH40 U50 ( .A1(wb_addr_o[27]), .A2(n36), .B1(cpu_addr_i[27]), .B2(
        n37), .Z(n120) );
  AO22V4_8TH40 U51 ( .A1(wb_addr_o[26]), .A2(n36), .B1(cpu_addr_i[26]), .B2(
        n37), .Z(n119) );
  AO22V4_8TH40 U52 ( .A1(wb_addr_o[25]), .A2(n36), .B1(cpu_addr_i[25]), .B2(
        n37), .Z(n118) );
  AO22V4_8TH40 U53 ( .A1(wb_addr_o[24]), .A2(n36), .B1(cpu_addr_i[24]), .B2(
        n37), .Z(n117) );
  AO22V4_8TH40 U54 ( .A1(wb_addr_o[23]), .A2(n36), .B1(cpu_addr_i[23]), .B2(
        n37), .Z(n116) );
  AO22V4_8TH40 U55 ( .A1(wb_addr_o[22]), .A2(n36), .B1(cpu_addr_i[22]), .B2(
        n37), .Z(n115) );
  AO22V4_8TH40 U56 ( .A1(wb_addr_o[21]), .A2(n36), .B1(cpu_addr_i[21]), .B2(
        n37), .Z(n114) );
  AO22V4_8TH40 U57 ( .A1(wb_addr_o[20]), .A2(n36), .B1(cpu_addr_i[20]), .B2(
        n37), .Z(n113) );
  AO22V4_8TH40 U58 ( .A1(wb_addr_o[19]), .A2(n36), .B1(cpu_addr_i[19]), .B2(
        n37), .Z(n112) );
  AO22V4_8TH40 U59 ( .A1(wb_addr_o[18]), .A2(n36), .B1(cpu_addr_i[18]), .B2(
        n37), .Z(n111) );
  AO22V4_8TH40 U60 ( .A1(wb_addr_o[17]), .A2(n36), .B1(cpu_addr_i[17]), .B2(
        n37), .Z(n110) );
  AO22V4_8TH40 U61 ( .A1(wb_addr_o[16]), .A2(n36), .B1(cpu_addr_i[16]), .B2(
        n37), .Z(n109) );
  AO22V4_8TH40 U62 ( .A1(wb_addr_o[15]), .A2(n36), .B1(cpu_addr_i[15]), .B2(
        n37), .Z(n108) );
  AO22V4_8TH40 U63 ( .A1(wb_addr_o[14]), .A2(n36), .B1(cpu_addr_i[14]), .B2(
        n37), .Z(n107) );
  AO22V4_8TH40 U64 ( .A1(wb_addr_o[13]), .A2(n36), .B1(cpu_addr_i[13]), .B2(
        n37), .Z(n106) );
  AO22V4_8TH40 U65 ( .A1(wb_addr_o[12]), .A2(n36), .B1(cpu_addr_i[12]), .B2(
        n37), .Z(n105) );
  AO22V4_8TH40 U66 ( .A1(wb_addr_o[11]), .A2(n36), .B1(cpu_addr_i[11]), .B2(
        n37), .Z(n104) );
  AO22V4_8TH40 U67 ( .A1(wb_addr_o[10]), .A2(n36), .B1(cpu_addr_i[10]), .B2(
        n37), .Z(n103) );
  AO22V4_8TH40 U68 ( .A1(wb_addr_o[9]), .A2(n36), .B1(cpu_addr_i[9]), .B2(n37), 
        .Z(n102) );
  AO22V4_8TH40 U69 ( .A1(wb_addr_o[8]), .A2(n36), .B1(cpu_addr_i[8]), .B2(n37), 
        .Z(n101) );
  AO22V4_8TH40 U70 ( .A1(wb_addr_o[7]), .A2(n36), .B1(cpu_addr_i[7]), .B2(n37), 
        .Z(n100) );
  INOR2V2_8TH40 U71 ( .A1(n86), .B1(n36), .ZN(n37) );
  OAI31V2_8TH40 U72 ( .A1(n43), .A2(n44), .A3(n41), .B(n36), .ZN(n40) );
  AO22V1_8TH40 U73 ( .A1(n36), .A2(wb_we_o), .B1(n37), .B2(cpu_we_i), .Z(n129)
         );
  NAND2V2_8TH40 U74 ( .A1(n38), .A2(n39), .ZN(n195) );
  AO33V0_8TH40 U75 ( .A1(n1), .A2(n2), .A3(n35), .B1(flush_i_BAR), .B2(n86), 
        .B3(cpu_ce_i), .Z(stall_req) );
  CLKNV1_8TH40 U76 ( .I(wb_ack_i), .ZN(n2) );
  MUX2NV0_8TH40 U77 ( .I0(wb_state[0]), .I1(n86), .S(n40), .ZN(n38) );
  OAI21V0_8TH40 U78 ( .A1(n41), .A2(n40), .B(n39), .ZN(n194) );
  OAI31V0_8TH40 U79 ( .A1(stall_ctrl[1]), .A2(stall_ctrl[4]), .A3(
        stall_ctrl[3]), .B(n42), .ZN(n39) );
  OR3V0_8TH40 U80 ( .A1(stall_ctrl[3]), .A2(stall_ctrl[4]), .A3(stall_ctrl[1]), 
        .Z(n43) );
  OAI22V0_8TH40 U81 ( .A1(n34), .A2(n45), .B1(n46), .B2(n47), .ZN(n193) );
  OAI22V0_8TH40 U82 ( .A1(n33), .A2(n45), .B1(n46), .B2(n48), .ZN(n192) );
  OAI22V0_8TH40 U83 ( .A1(n32), .A2(n45), .B1(n46), .B2(n49), .ZN(n191) );
  OAI22V0_8TH40 U84 ( .A1(n31), .A2(n45), .B1(n46), .B2(n50), .ZN(n190) );
  OAI22V0_8TH40 U85 ( .A1(n30), .A2(n45), .B1(n46), .B2(n51), .ZN(n189) );
  OAI22V0_8TH40 U86 ( .A1(n29), .A2(n45), .B1(n46), .B2(n52), .ZN(n188) );
  OAI22V0_8TH40 U87 ( .A1(n28), .A2(n45), .B1(n46), .B2(n53), .ZN(n187) );
  OAI22V0_8TH40 U88 ( .A1(n27), .A2(n45), .B1(n46), .B2(n54), .ZN(n186) );
  OAI22V0_8TH40 U89 ( .A1(n26), .A2(n45), .B1(n46), .B2(n55), .ZN(n185) );
  OAI22V0_8TH40 U90 ( .A1(n25), .A2(n45), .B1(n46), .B2(n56), .ZN(n184) );
  OAI22V0_8TH40 U91 ( .A1(n24), .A2(n45), .B1(n46), .B2(n57), .ZN(n183) );
  OAI22V0_8TH40 U92 ( .A1(n23), .A2(n45), .B1(n46), .B2(n58), .ZN(n182) );
  OAI22V0_8TH40 U93 ( .A1(n22), .A2(n45), .B1(n46), .B2(n59), .ZN(n181) );
  OAI22V0_8TH40 U94 ( .A1(n21), .A2(n45), .B1(n46), .B2(n60), .ZN(n180) );
  OAI22V0_8TH40 U95 ( .A1(n20), .A2(n45), .B1(n46), .B2(n61), .ZN(n179) );
  OAI22V0_8TH40 U96 ( .A1(n19), .A2(n45), .B1(n46), .B2(n62), .ZN(n178) );
  OAI22V0_8TH40 U97 ( .A1(n18), .A2(n45), .B1(n46), .B2(n63), .ZN(n177) );
  OAI22V0_8TH40 U98 ( .A1(n17), .A2(n45), .B1(n46), .B2(n64), .ZN(n176) );
  OAI22V0_8TH40 U99 ( .A1(n16), .A2(n45), .B1(n46), .B2(n65), .ZN(n175) );
  OAI22V0_8TH40 U100 ( .A1(n15), .A2(n45), .B1(n46), .B2(n66), .ZN(n174) );
  OAI22V0_8TH40 U101 ( .A1(n14), .A2(n45), .B1(n46), .B2(n67), .ZN(n173) );
  OAI22V0_8TH40 U102 ( .A1(n13), .A2(n45), .B1(n46), .B2(n68), .ZN(n172) );
  OAI22V0_8TH40 U103 ( .A1(n12), .A2(n45), .B1(n46), .B2(n69), .ZN(n171) );
  OAI22V0_8TH40 U104 ( .A1(n11), .A2(n45), .B1(n46), .B2(n70), .ZN(n170) );
  OAI22V0_8TH40 U105 ( .A1(n10), .A2(n45), .B1(n46), .B2(n71), .ZN(n169) );
  OAI22V0_8TH40 U106 ( .A1(n9), .A2(n45), .B1(n46), .B2(n72), .ZN(n168) );
  OAI22V0_8TH40 U107 ( .A1(n8), .A2(n45), .B1(n46), .B2(n73), .ZN(n167) );
  OAI22V0_8TH40 U108 ( .A1(n7), .A2(n45), .B1(n46), .B2(n74), .ZN(n166) );
  OAI22V0_8TH40 U109 ( .A1(n6), .A2(n45), .B1(n46), .B2(n75), .ZN(n165) );
  OAI22V0_8TH40 U110 ( .A1(n5), .A2(n45), .B1(n46), .B2(n76), .ZN(n164) );
  OAI22V0_8TH40 U111 ( .A1(n4), .A2(n45), .B1(n46), .B2(n77), .ZN(n163) );
  OAI22V0_8TH40 U112 ( .A1(n3), .A2(n45), .B1(n46), .B2(n78), .ZN(n162) );
  CLKNAND2V1_8TH40 U113 ( .A1(n42), .A2(n45), .ZN(n46) );
  OAI221V0_8TH40 U114 ( .A1(wb_ack_i), .A2(n79), .B1(cpu_we_i), .B2(n80), .C(
        n81), .ZN(n45) );
  NOR3V0P5_8TH40 U115 ( .A1(wb_state[0]), .A2(wb_state[1]), .A3(rst), .ZN(n86)
         );
  CLKNV1_8TH40 U116 ( .I(n85), .ZN(n36) );
  NAND3V0P5_8TH40 U117 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n85) );
  INAND2V0_8TH40 U118 ( .A1(flush_i_BAR), .B1(n1), .ZN(n79) );
  OAI22V0_8TH40 U119 ( .A1(n78), .A2(n82), .B1(n3), .B2(n83), .ZN(N419) );
  CLKNV1_8TH40 U120 ( .I(wb_data_i[31]), .ZN(n78) );
  OAI22V0_8TH40 U121 ( .A1(n77), .A2(n82), .B1(n4), .B2(n83), .ZN(N418) );
  CLKNV1_8TH40 U122 ( .I(wb_data_i[30]), .ZN(n77) );
  OAI22V0_8TH40 U123 ( .A1(n76), .A2(n82), .B1(n5), .B2(n83), .ZN(N417) );
  CLKNV1_8TH40 U124 ( .I(wb_data_i[29]), .ZN(n76) );
  OAI22V0_8TH40 U125 ( .A1(n75), .A2(n82), .B1(n6), .B2(n83), .ZN(N416) );
  CLKNV1_8TH40 U126 ( .I(wb_data_i[28]), .ZN(n75) );
  OAI22V0_8TH40 U127 ( .A1(n74), .A2(n82), .B1(n7), .B2(n83), .ZN(N415) );
  CLKNV1_8TH40 U128 ( .I(wb_data_i[27]), .ZN(n74) );
  OAI22V0_8TH40 U129 ( .A1(n73), .A2(n82), .B1(n8), .B2(n83), .ZN(N414) );
  CLKNV1_8TH40 U130 ( .I(wb_data_i[26]), .ZN(n73) );
  OAI22V0_8TH40 U131 ( .A1(n72), .A2(n82), .B1(n9), .B2(n83), .ZN(N413) );
  CLKNV1_8TH40 U132 ( .I(wb_data_i[25]), .ZN(n72) );
  OAI22V0_8TH40 U133 ( .A1(n71), .A2(n82), .B1(n10), .B2(n83), .ZN(N412) );
  CLKNV1_8TH40 U134 ( .I(wb_data_i[24]), .ZN(n71) );
  OAI22V0_8TH40 U135 ( .A1(n70), .A2(n82), .B1(n11), .B2(n83), .ZN(N411) );
  CLKNV1_8TH40 U136 ( .I(wb_data_i[23]), .ZN(n70) );
  OAI22V0_8TH40 U137 ( .A1(n69), .A2(n82), .B1(n12), .B2(n83), .ZN(N410) );
  CLKNV1_8TH40 U138 ( .I(wb_data_i[22]), .ZN(n69) );
  OAI22V0_8TH40 U139 ( .A1(n68), .A2(n82), .B1(n13), .B2(n83), .ZN(N409) );
  CLKNV1_8TH40 U140 ( .I(wb_data_i[21]), .ZN(n68) );
  OAI22V0_8TH40 U141 ( .A1(n67), .A2(n82), .B1(n14), .B2(n83), .ZN(N408) );
  CLKNV1_8TH40 U142 ( .I(wb_data_i[20]), .ZN(n67) );
  OAI22V0_8TH40 U143 ( .A1(n66), .A2(n82), .B1(n15), .B2(n83), .ZN(N407) );
  CLKNV1_8TH40 U144 ( .I(wb_data_i[19]), .ZN(n66) );
  OAI22V0_8TH40 U145 ( .A1(n65), .A2(n82), .B1(n16), .B2(n83), .ZN(N406) );
  CLKNV1_8TH40 U146 ( .I(wb_data_i[18]), .ZN(n65) );
  OAI22V0_8TH40 U147 ( .A1(n64), .A2(n82), .B1(n17), .B2(n83), .ZN(N405) );
  CLKNV1_8TH40 U148 ( .I(wb_data_i[17]), .ZN(n64) );
  OAI22V0_8TH40 U149 ( .A1(n63), .A2(n82), .B1(n18), .B2(n83), .ZN(N404) );
  CLKNV1_8TH40 U150 ( .I(wb_data_i[16]), .ZN(n63) );
  OAI22V0_8TH40 U151 ( .A1(n62), .A2(n82), .B1(n19), .B2(n83), .ZN(N403) );
  CLKNV1_8TH40 U152 ( .I(wb_data_i[15]), .ZN(n62) );
  OAI22V0_8TH40 U153 ( .A1(n61), .A2(n82), .B1(n20), .B2(n83), .ZN(N402) );
  CLKNV1_8TH40 U154 ( .I(wb_data_i[14]), .ZN(n61) );
  OAI22V0_8TH40 U155 ( .A1(n60), .A2(n82), .B1(n21), .B2(n83), .ZN(N401) );
  CLKNV1_8TH40 U156 ( .I(wb_data_i[13]), .ZN(n60) );
  OAI22V0_8TH40 U157 ( .A1(n59), .A2(n82), .B1(n22), .B2(n83), .ZN(N400) );
  CLKNV1_8TH40 U158 ( .I(wb_data_i[12]), .ZN(n59) );
  OAI22V0_8TH40 U159 ( .A1(n58), .A2(n82), .B1(n23), .B2(n83), .ZN(N399) );
  CLKNV1_8TH40 U160 ( .I(wb_data_i[11]), .ZN(n58) );
  OAI22V0_8TH40 U161 ( .A1(n57), .A2(n82), .B1(n24), .B2(n83), .ZN(N398) );
  CLKNV1_8TH40 U162 ( .I(wb_data_i[10]), .ZN(n57) );
  OAI22V0_8TH40 U163 ( .A1(n56), .A2(n82), .B1(n25), .B2(n83), .ZN(N397) );
  CLKNV1_8TH40 U164 ( .I(wb_data_i[9]), .ZN(n56) );
  OAI22V0_8TH40 U165 ( .A1(n55), .A2(n82), .B1(n26), .B2(n83), .ZN(N396) );
  CLKNV1_8TH40 U166 ( .I(wb_data_i[8]), .ZN(n55) );
  OAI22V0_8TH40 U167 ( .A1(n54), .A2(n82), .B1(n27), .B2(n83), .ZN(N395) );
  CLKNV1_8TH40 U168 ( .I(wb_data_i[7]), .ZN(n54) );
  OAI22V0_8TH40 U169 ( .A1(n53), .A2(n82), .B1(n28), .B2(n83), .ZN(N394) );
  CLKNV1_8TH40 U170 ( .I(wb_data_i[6]), .ZN(n53) );
  OAI22V0_8TH40 U171 ( .A1(n52), .A2(n82), .B1(n29), .B2(n83), .ZN(N393) );
  CLKNV1_8TH40 U172 ( .I(wb_data_i[5]), .ZN(n52) );
  OAI22V0_8TH40 U173 ( .A1(n51), .A2(n82), .B1(n30), .B2(n83), .ZN(N392) );
  CLKNV1_8TH40 U174 ( .I(wb_data_i[4]), .ZN(n51) );
  OAI22V0_8TH40 U175 ( .A1(n50), .A2(n82), .B1(n31), .B2(n83), .ZN(N391) );
  CLKNV1_8TH40 U176 ( .I(wb_data_i[3]), .ZN(n50) );
  OAI22V0_8TH40 U177 ( .A1(n49), .A2(n82), .B1(n32), .B2(n83), .ZN(N390) );
  CLKNV1_8TH40 U178 ( .I(wb_data_i[2]), .ZN(n49) );
  OAI22V0_8TH40 U179 ( .A1(n48), .A2(n82), .B1(n33), .B2(n83), .ZN(N389) );
  CLKNV1_8TH40 U180 ( .I(wb_data_i[1]), .ZN(n48) );
  OAI22V0_8TH40 U181 ( .A1(n47), .A2(n82), .B1(n34), .B2(n83), .ZN(N388) );
  NAND3V0P5_8TH40 U182 ( .A1(wb_state[0]), .A2(n35), .A3(wb_state[1]), .ZN(n83) );
  INAND2V0_8TH40 U183 ( .A1(wb_we_o), .B1(n42), .ZN(n82) );
  NOR2V0P5_8TH40 U184 ( .A1(n80), .A2(rst), .ZN(n42) );
  CLKNAND2V1_8TH40 U185 ( .A1(wb_ack_i), .A2(n1), .ZN(n80) );
  NOR2V0P5_8TH40 U186 ( .A1(n44), .A2(wb_state[1]), .ZN(n1) );
  CLKNV1_8TH40 U187 ( .I(wb_data_i[0]), .ZN(n47) );
  CLKNAND2V1_8TH40 U188 ( .A1(n81), .A2(n44), .ZN(N387) );
  AND2V0_8TH40 U189 ( .A1(n84), .A2(n35), .Z(n81) );
  CLKNV1_8TH40 U190 ( .I(rst), .ZN(n35) );
  NAND4V0P5_8TH40 U191 ( .A1(flush_i_BAR), .A2(cpu_ce_i), .A3(n44), .A4(n41), 
        .ZN(n84) );
  CLKNV1_8TH40 U192 ( .I(wb_state[1]), .ZN(n41) );
  CLKNV1_8TH40 U193 ( .I(wb_state[0]), .ZN(n44) );
endmodule


module wb_interface_1 ( clk, rst, stall_ctrl, cpu_ce_i, cpu_data_i, cpu_addr_i, 
        cpu_we_i, cpu_sel_i, cpu_data_o, wb_data_i, wb_ack_i, wb_addr_o, 
        wb_data_o, wb_we_o, wb_sel_o, wb_stb_o, wb_cyc_o, stall_req, 
        flush_i_BAR );
  input [5:0] stall_ctrl;
  input [31:0] cpu_data_i;
  input [31:0] cpu_addr_i;
  input [3:0] cpu_sel_i;
  output [31:0] cpu_data_o;
  input [31:0] wb_data_i;
  output [31:0] wb_addr_o;
  output [31:0] wb_data_o;
  output [3:0] wb_sel_o;
  input clk, rst, cpu_ce_i, cpu_we_i, wb_ack_i, flush_i_BAR;
  output wb_we_o, wb_stb_o, wb_cyc_o, stall_req;
  wire   N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, n1,
         n2, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287;
  wire   [1:0] wb_state;

  DQV4_8TH40 wb_state_reg_0_ ( .D(n157), .CK(clk), .Q(wb_state[0]) );
  DQV4_8TH40 wb_state_reg_1_ ( .D(n158), .CK(clk), .Q(wb_state[1]) );
  DQNV4_8TH40 data_buf_reg_31_ ( .D(n219), .CK(clk), .QN(n287) );
  DQNV4_8TH40 data_buf_reg_30_ ( .D(n218), .CK(clk), .QN(n286) );
  DQNV4_8TH40 data_buf_reg_29_ ( .D(n217), .CK(clk), .QN(n285) );
  DQNV4_8TH40 data_buf_reg_28_ ( .D(n216), .CK(clk), .QN(n284) );
  DQNV4_8TH40 data_buf_reg_27_ ( .D(n215), .CK(clk), .QN(n283) );
  DQNV4_8TH40 data_buf_reg_26_ ( .D(n214), .CK(clk), .QN(n282) );
  DQNV4_8TH40 data_buf_reg_25_ ( .D(n213), .CK(clk), .QN(n281) );
  DQNV4_8TH40 data_buf_reg_24_ ( .D(n212), .CK(clk), .QN(n280) );
  DQNV4_8TH40 data_buf_reg_23_ ( .D(n211), .CK(clk), .QN(n279) );
  DQNV4_8TH40 data_buf_reg_22_ ( .D(n210), .CK(clk), .QN(n278) );
  DQNV4_8TH40 data_buf_reg_21_ ( .D(n209), .CK(clk), .QN(n277) );
  DQNV4_8TH40 data_buf_reg_20_ ( .D(n208), .CK(clk), .QN(n276) );
  DQNV4_8TH40 data_buf_reg_19_ ( .D(n207), .CK(clk), .QN(n275) );
  DQNV4_8TH40 data_buf_reg_18_ ( .D(n206), .CK(clk), .QN(n274) );
  DQNV4_8TH40 data_buf_reg_17_ ( .D(n205), .CK(clk), .QN(n273) );
  DQNV4_8TH40 data_buf_reg_16_ ( .D(n204), .CK(clk), .QN(n272) );
  DQNV4_8TH40 data_buf_reg_15_ ( .D(n203), .CK(clk), .QN(n271) );
  DQNV4_8TH40 data_buf_reg_14_ ( .D(n202), .CK(clk), .QN(n270) );
  DQNV4_8TH40 data_buf_reg_13_ ( .D(n201), .CK(clk), .QN(n269) );
  DQNV4_8TH40 data_buf_reg_12_ ( .D(n200), .CK(clk), .QN(n268) );
  DQNV4_8TH40 data_buf_reg_11_ ( .D(n199), .CK(clk), .QN(n267) );
  DQNV4_8TH40 data_buf_reg_10_ ( .D(n198), .CK(clk), .QN(n266) );
  DQNV4_8TH40 data_buf_reg_9_ ( .D(n197), .CK(clk), .QN(n265) );
  DQNV4_8TH40 data_buf_reg_8_ ( .D(n196), .CK(clk), .QN(n264) );
  DQNV4_8TH40 data_buf_reg_7_ ( .D(n195), .CK(clk), .QN(n263) );
  DQNV4_8TH40 data_buf_reg_6_ ( .D(n194), .CK(clk), .QN(n262) );
  DQNV4_8TH40 data_buf_reg_5_ ( .D(n193), .CK(clk), .QN(n261) );
  DQNV4_8TH40 data_buf_reg_4_ ( .D(n192), .CK(clk), .QN(n260) );
  DQNV4_8TH40 data_buf_reg_3_ ( .D(n191), .CK(clk), .QN(n259) );
  DQNV4_8TH40 data_buf_reg_2_ ( .D(n161), .CK(clk), .QN(n258) );
  DQNV4_8TH40 data_buf_reg_1_ ( .D(n160), .CK(clk), .QN(n257) );
  DQNV4_8TH40 data_buf_reg_0_ ( .D(n159), .CK(clk), .QN(n256) );
  DQV4_8TH40 wb_sel_o_reg_3_ ( .D(n223), .CK(clk), .Q(wb_sel_o[3]) );
  DQV4_8TH40 wb_sel_o_reg_2_ ( .D(n222), .CK(clk), .Q(wb_sel_o[2]) );
  DQV4_8TH40 wb_sel_o_reg_1_ ( .D(n221), .CK(clk), .Q(wb_sel_o[1]) );
  DQV4_8TH40 wb_sel_o_reg_0_ ( .D(n220), .CK(clk), .Q(wb_sel_o[0]) );
  DQV4_8TH40 wb_we_o_reg ( .D(n86), .CK(clk), .Q(wb_we_o) );
  DQV4_8TH40 wb_data_o_reg_31_ ( .D(n154), .CK(clk), .Q(wb_data_o[31]) );
  DQV4_8TH40 wb_data_o_reg_30_ ( .D(n153), .CK(clk), .Q(wb_data_o[30]) );
  DQV4_8TH40 wb_data_o_reg_29_ ( .D(n152), .CK(clk), .Q(wb_data_o[29]) );
  DQV4_8TH40 wb_data_o_reg_28_ ( .D(n151), .CK(clk), .Q(wb_data_o[28]) );
  DQV4_8TH40 wb_data_o_reg_27_ ( .D(n150), .CK(clk), .Q(wb_data_o[27]) );
  DQV4_8TH40 wb_data_o_reg_26_ ( .D(n149), .CK(clk), .Q(wb_data_o[26]) );
  DQV4_8TH40 wb_data_o_reg_25_ ( .D(n148), .CK(clk), .Q(wb_data_o[25]) );
  DQV4_8TH40 wb_data_o_reg_24_ ( .D(n147), .CK(clk), .Q(wb_data_o[24]) );
  DQV4_8TH40 wb_data_o_reg_23_ ( .D(n146), .CK(clk), .Q(wb_data_o[23]) );
  DQV4_8TH40 wb_data_o_reg_22_ ( .D(n145), .CK(clk), .Q(wb_data_o[22]) );
  DQV4_8TH40 wb_data_o_reg_21_ ( .D(n144), .CK(clk), .Q(wb_data_o[21]) );
  DQV4_8TH40 wb_data_o_reg_20_ ( .D(n143), .CK(clk), .Q(wb_data_o[20]) );
  DQV4_8TH40 wb_data_o_reg_19_ ( .D(n142), .CK(clk), .Q(wb_data_o[19]) );
  DQV4_8TH40 wb_data_o_reg_18_ ( .D(n141), .CK(clk), .Q(wb_data_o[18]) );
  DQV4_8TH40 wb_data_o_reg_17_ ( .D(n140), .CK(clk), .Q(wb_data_o[17]) );
  DQV4_8TH40 wb_data_o_reg_16_ ( .D(n139), .CK(clk), .Q(wb_data_o[16]) );
  DQV4_8TH40 wb_data_o_reg_15_ ( .D(n138), .CK(clk), .Q(wb_data_o[15]) );
  DQV4_8TH40 wb_data_o_reg_14_ ( .D(n137), .CK(clk), .Q(wb_data_o[14]) );
  DQV4_8TH40 wb_data_o_reg_13_ ( .D(n136), .CK(clk), .Q(wb_data_o[13]) );
  DQV4_8TH40 wb_data_o_reg_12_ ( .D(n135), .CK(clk), .Q(wb_data_o[12]) );
  DQV4_8TH40 wb_data_o_reg_11_ ( .D(n134), .CK(clk), .Q(wb_data_o[11]) );
  DQV4_8TH40 wb_data_o_reg_10_ ( .D(n133), .CK(clk), .Q(wb_data_o[10]) );
  DQV4_8TH40 wb_data_o_reg_9_ ( .D(n132), .CK(clk), .Q(wb_data_o[9]) );
  DQV4_8TH40 wb_data_o_reg_8_ ( .D(n131), .CK(clk), .Q(wb_data_o[8]) );
  DQV4_8TH40 wb_data_o_reg_7_ ( .D(n130), .CK(clk), .Q(wb_data_o[7]) );
  DQV4_8TH40 wb_data_o_reg_6_ ( .D(n129), .CK(clk), .Q(wb_data_o[6]) );
  DQV4_8TH40 wb_data_o_reg_5_ ( .D(n92), .CK(clk), .Q(wb_data_o[5]) );
  DQV4_8TH40 wb_data_o_reg_4_ ( .D(n91), .CK(clk), .Q(wb_data_o[4]) );
  DQV4_8TH40 wb_data_o_reg_3_ ( .D(n90), .CK(clk), .Q(wb_data_o[3]) );
  DQV4_8TH40 wb_data_o_reg_2_ ( .D(n89), .CK(clk), .Q(wb_data_o[2]) );
  DQV4_8TH40 wb_data_o_reg_1_ ( .D(n88), .CK(clk), .Q(wb_data_o[1]) );
  DQV4_8TH40 wb_data_o_reg_0_ ( .D(n87), .CK(clk), .Q(wb_data_o[0]) );
  DQV4_8TH40 wb_addr_o_reg_31_ ( .D(n224), .CK(clk), .Q(wb_addr_o[31]) );
  DQV4_8TH40 wb_addr_o_reg_30_ ( .D(n225), .CK(clk), .Q(wb_addr_o[30]) );
  DQV4_8TH40 wb_addr_o_reg_29_ ( .D(n226), .CK(clk), .Q(wb_addr_o[29]) );
  DQV4_8TH40 wb_addr_o_reg_28_ ( .D(n227), .CK(clk), .Q(wb_addr_o[28]) );
  DQV4_8TH40 wb_addr_o_reg_27_ ( .D(n228), .CK(clk), .Q(wb_addr_o[27]) );
  DQV4_8TH40 wb_addr_o_reg_26_ ( .D(n229), .CK(clk), .Q(wb_addr_o[26]) );
  DQV4_8TH40 wb_addr_o_reg_25_ ( .D(n230), .CK(clk), .Q(wb_addr_o[25]) );
  DQV4_8TH40 wb_addr_o_reg_24_ ( .D(n231), .CK(clk), .Q(wb_addr_o[24]) );
  DQV4_8TH40 wb_addr_o_reg_23_ ( .D(n232), .CK(clk), .Q(wb_addr_o[23]) );
  DQV4_8TH40 wb_addr_o_reg_22_ ( .D(n233), .CK(clk), .Q(wb_addr_o[22]) );
  DQV4_8TH40 wb_addr_o_reg_21_ ( .D(n234), .CK(clk), .Q(wb_addr_o[21]) );
  DQV4_8TH40 wb_addr_o_reg_20_ ( .D(n235), .CK(clk), .Q(wb_addr_o[20]) );
  DQV4_8TH40 wb_addr_o_reg_19_ ( .D(n236), .CK(clk), .Q(wb_addr_o[19]) );
  DQV4_8TH40 wb_addr_o_reg_18_ ( .D(n237), .CK(clk), .Q(wb_addr_o[18]) );
  DQV4_8TH40 wb_addr_o_reg_17_ ( .D(n238), .CK(clk), .Q(wb_addr_o[17]) );
  DQV4_8TH40 wb_addr_o_reg_16_ ( .D(n239), .CK(clk), .Q(wb_addr_o[16]) );
  DQV4_8TH40 wb_addr_o_reg_15_ ( .D(n240), .CK(clk), .Q(wb_addr_o[15]) );
  DQV4_8TH40 wb_addr_o_reg_14_ ( .D(n241), .CK(clk), .Q(wb_addr_o[14]) );
  DQV4_8TH40 wb_addr_o_reg_13_ ( .D(n242), .CK(clk), .Q(wb_addr_o[13]) );
  DQV4_8TH40 wb_addr_o_reg_12_ ( .D(n243), .CK(clk), .Q(wb_addr_o[12]) );
  DQV4_8TH40 wb_addr_o_reg_11_ ( .D(n244), .CK(clk), .Q(wb_addr_o[11]) );
  DQV4_8TH40 wb_addr_o_reg_10_ ( .D(n245), .CK(clk), .Q(wb_addr_o[10]) );
  DQV4_8TH40 wb_addr_o_reg_9_ ( .D(n246), .CK(clk), .Q(wb_addr_o[9]) );
  DQV4_8TH40 wb_addr_o_reg_8_ ( .D(n247), .CK(clk), .Q(wb_addr_o[8]) );
  DQV4_8TH40 wb_addr_o_reg_7_ ( .D(n248), .CK(clk), .Q(wb_addr_o[7]) );
  DQV4_8TH40 wb_addr_o_reg_6_ ( .D(n249), .CK(clk), .Q(wb_addr_o[6]) );
  DQV4_8TH40 wb_addr_o_reg_5_ ( .D(n250), .CK(clk), .Q(wb_addr_o[5]) );
  DQV4_8TH40 wb_addr_o_reg_4_ ( .D(n251), .CK(clk), .Q(wb_addr_o[4]) );
  DQV4_8TH40 wb_addr_o_reg_3_ ( .D(n252), .CK(clk), .Q(wb_addr_o[3]) );
  DQV4_8TH40 wb_addr_o_reg_2_ ( .D(n253), .CK(clk), .Q(wb_addr_o[2]) );
  DQV4_8TH40 wb_addr_o_reg_1_ ( .D(n254), .CK(clk), .Q(wb_addr_o[1]) );
  DQV4_8TH40 wb_addr_o_reg_0_ ( .D(n255), .CK(clk), .Q(wb_addr_o[0]) );
  EDQV2_8TH40 wb_cyc_o_reg ( .D(n156), .E(n155), .CK(clk), .Q(wb_cyc_o) );
  EDQV2_8TH40 wb_stb_o_reg ( .D(n156), .E(n155), .CK(clk), .Q(wb_stb_o) );
  LAHQV4_8TH40 cpu_data_o_reg_31_ ( .E(N387), .D(N419), .Q(cpu_data_o[31]) );
  LAHQV4_8TH40 cpu_data_o_reg_30_ ( .E(N387), .D(N418), .Q(cpu_data_o[30]) );
  LAHQV4_8TH40 cpu_data_o_reg_29_ ( .E(N387), .D(N417), .Q(cpu_data_o[29]) );
  LAHQV4_8TH40 cpu_data_o_reg_28_ ( .E(N387), .D(N416), .Q(cpu_data_o[28]) );
  LAHQV4_8TH40 cpu_data_o_reg_27_ ( .E(N387), .D(N415), .Q(cpu_data_o[27]) );
  LAHQV4_8TH40 cpu_data_o_reg_26_ ( .E(N387), .D(N414), .Q(cpu_data_o[26]) );
  LAHQV4_8TH40 cpu_data_o_reg_25_ ( .E(N387), .D(N413), .Q(cpu_data_o[25]) );
  LAHQV4_8TH40 cpu_data_o_reg_24_ ( .E(N387), .D(N412), .Q(cpu_data_o[24]) );
  LAHQV4_8TH40 cpu_data_o_reg_23_ ( .E(N387), .D(N411), .Q(cpu_data_o[23]) );
  LAHQV4_8TH40 cpu_data_o_reg_22_ ( .E(N387), .D(N410), .Q(cpu_data_o[22]) );
  LAHQV4_8TH40 cpu_data_o_reg_21_ ( .E(N387), .D(N409), .Q(cpu_data_o[21]) );
  LAHQV4_8TH40 cpu_data_o_reg_20_ ( .E(N387), .D(N408), .Q(cpu_data_o[20]) );
  LAHQV4_8TH40 cpu_data_o_reg_19_ ( .E(N387), .D(N407), .Q(cpu_data_o[19]) );
  LAHQV4_8TH40 cpu_data_o_reg_18_ ( .E(N387), .D(N406), .Q(cpu_data_o[18]) );
  LAHQV4_8TH40 cpu_data_o_reg_17_ ( .E(N387), .D(N405), .Q(cpu_data_o[17]) );
  LAHQV4_8TH40 cpu_data_o_reg_16_ ( .E(N387), .D(N404), .Q(cpu_data_o[16]) );
  LAHQV4_8TH40 cpu_data_o_reg_15_ ( .E(N387), .D(N403), .Q(cpu_data_o[15]) );
  LAHQV4_8TH40 cpu_data_o_reg_14_ ( .E(N387), .D(N402), .Q(cpu_data_o[14]) );
  LAHQV4_8TH40 cpu_data_o_reg_13_ ( .E(N387), .D(N401), .Q(cpu_data_o[13]) );
  LAHQV4_8TH40 cpu_data_o_reg_12_ ( .E(N387), .D(N400), .Q(cpu_data_o[12]) );
  LAHQV4_8TH40 cpu_data_o_reg_11_ ( .E(N387), .D(N399), .Q(cpu_data_o[11]) );
  LAHQV4_8TH40 cpu_data_o_reg_10_ ( .E(N387), .D(N398), .Q(cpu_data_o[10]) );
  LAHQV4_8TH40 cpu_data_o_reg_9_ ( .E(N387), .D(N397), .Q(cpu_data_o[9]) );
  LAHQV4_8TH40 cpu_data_o_reg_8_ ( .E(N387), .D(N396), .Q(cpu_data_o[8]) );
  LAHQV4_8TH40 cpu_data_o_reg_7_ ( .E(N387), .D(N395), .Q(cpu_data_o[7]) );
  LAHQV4_8TH40 cpu_data_o_reg_6_ ( .E(N387), .D(N394), .Q(cpu_data_o[6]) );
  LAHQV4_8TH40 cpu_data_o_reg_5_ ( .E(N387), .D(N393), .Q(cpu_data_o[5]) );
  LAHQV4_8TH40 cpu_data_o_reg_4_ ( .E(N387), .D(N392), .Q(cpu_data_o[4]) );
  LAHQV4_8TH40 cpu_data_o_reg_3_ ( .E(N387), .D(N391), .Q(cpu_data_o[3]) );
  LAHQV4_8TH40 cpu_data_o_reg_2_ ( .E(N387), .D(N390), .Q(cpu_data_o[2]) );
  LAHQV4_8TH40 cpu_data_o_reg_1_ ( .E(N387), .D(N389), .Q(cpu_data_o[1]) );
  LAHQV4_8TH40 cpu_data_o_reg_0_ ( .E(N387), .D(N388), .Q(cpu_data_o[0]) );
  AO22V4_8TH40 U3 ( .A1(wb_addr_o[0]), .A2(n37), .B1(cpu_addr_i[0]), .B2(n38), 
        .Z(n255) );
  AO22V4_8TH40 U4 ( .A1(wb_addr_o[1]), .A2(n37), .B1(cpu_addr_i[1]), .B2(n38), 
        .Z(n254) );
  AO22V4_8TH40 U5 ( .A1(wb_addr_o[2]), .A2(n37), .B1(cpu_addr_i[2]), .B2(n38), 
        .Z(n253) );
  AO22V4_8TH40 U6 ( .A1(wb_addr_o[3]), .A2(n37), .B1(cpu_addr_i[3]), .B2(n38), 
        .Z(n252) );
  AO22V4_8TH40 U7 ( .A1(wb_addr_o[4]), .A2(n37), .B1(cpu_addr_i[4]), .B2(n38), 
        .Z(n251) );
  AO22V4_8TH40 U8 ( .A1(wb_addr_o[5]), .A2(n37), .B1(cpu_addr_i[5]), .B2(n38), 
        .Z(n250) );
  AO22V4_8TH40 U9 ( .A1(wb_addr_o[6]), .A2(n37), .B1(cpu_addr_i[6]), .B2(n38), 
        .Z(n249) );
  AO22V4_8TH40 U10 ( .A1(wb_addr_o[7]), .A2(n37), .B1(cpu_addr_i[7]), .B2(n38), 
        .Z(n248) );
  AO22V4_8TH40 U11 ( .A1(wb_addr_o[8]), .A2(n37), .B1(cpu_addr_i[8]), .B2(n38), 
        .Z(n247) );
  AO22V4_8TH40 U12 ( .A1(wb_addr_o[9]), .A2(n37), .B1(cpu_addr_i[9]), .B2(n38), 
        .Z(n246) );
  AO22V4_8TH40 U13 ( .A1(wb_addr_o[10]), .A2(n37), .B1(cpu_addr_i[10]), .B2(
        n38), .Z(n245) );
  AO22V4_8TH40 U14 ( .A1(wb_addr_o[11]), .A2(n37), .B1(cpu_addr_i[11]), .B2(
        n38), .Z(n244) );
  AO22V4_8TH40 U15 ( .A1(wb_addr_o[12]), .A2(n37), .B1(cpu_addr_i[12]), .B2(
        n38), .Z(n243) );
  AO22V4_8TH40 U16 ( .A1(wb_addr_o[13]), .A2(n37), .B1(cpu_addr_i[13]), .B2(
        n38), .Z(n242) );
  AO22V4_8TH40 U17 ( .A1(wb_addr_o[14]), .A2(n37), .B1(cpu_addr_i[14]), .B2(
        n38), .Z(n241) );
  AO22V4_8TH40 U18 ( .A1(wb_addr_o[15]), .A2(n37), .B1(cpu_addr_i[15]), .B2(
        n38), .Z(n240) );
  AO22V4_8TH40 U19 ( .A1(wb_addr_o[16]), .A2(n37), .B1(cpu_addr_i[16]), .B2(
        n38), .Z(n239) );
  AO22V4_8TH40 U20 ( .A1(wb_addr_o[17]), .A2(n37), .B1(cpu_addr_i[17]), .B2(
        n38), .Z(n238) );
  AO22V4_8TH40 U21 ( .A1(wb_addr_o[18]), .A2(n37), .B1(cpu_addr_i[18]), .B2(
        n38), .Z(n237) );
  AO22V4_8TH40 U22 ( .A1(wb_addr_o[19]), .A2(n37), .B1(cpu_addr_i[19]), .B2(
        n38), .Z(n236) );
  AO22V4_8TH40 U23 ( .A1(wb_addr_o[20]), .A2(n37), .B1(cpu_addr_i[20]), .B2(
        n38), .Z(n235) );
  AO22V4_8TH40 U24 ( .A1(wb_addr_o[21]), .A2(n37), .B1(cpu_addr_i[21]), .B2(
        n38), .Z(n234) );
  AO22V4_8TH40 U25 ( .A1(wb_addr_o[22]), .A2(n37), .B1(cpu_addr_i[22]), .B2(
        n38), .Z(n233) );
  AO22V4_8TH40 U26 ( .A1(wb_addr_o[23]), .A2(n37), .B1(cpu_addr_i[23]), .B2(
        n38), .Z(n232) );
  AO22V4_8TH40 U27 ( .A1(wb_addr_o[24]), .A2(n37), .B1(cpu_addr_i[24]), .B2(
        n38), .Z(n231) );
  AO22V4_8TH40 U28 ( .A1(wb_addr_o[25]), .A2(n37), .B1(cpu_addr_i[25]), .B2(
        n38), .Z(n230) );
  AO22V4_8TH40 U29 ( .A1(wb_addr_o[26]), .A2(n37), .B1(cpu_addr_i[26]), .B2(
        n38), .Z(n229) );
  AO22V4_8TH40 U30 ( .A1(wb_addr_o[27]), .A2(n37), .B1(cpu_addr_i[27]), .B2(
        n38), .Z(n228) );
  AO22V4_8TH40 U31 ( .A1(wb_addr_o[28]), .A2(n37), .B1(cpu_addr_i[28]), .B2(
        n38), .Z(n227) );
  AO22V4_8TH40 U32 ( .A1(wb_addr_o[29]), .A2(n37), .B1(cpu_addr_i[29]), .B2(
        n38), .Z(n226) );
  AO22V4_8TH40 U33 ( .A1(wb_addr_o[30]), .A2(n37), .B1(cpu_addr_i[30]), .B2(
        n38), .Z(n225) );
  AO22V4_8TH40 U34 ( .A1(wb_addr_o[31]), .A2(n37), .B1(cpu_addr_i[31]), .B2(
        n38), .Z(n224) );
  IOA21V8_8TH40 U35 ( .A1(wb_sel_o[0]), .A2(n37), .B(n79), .ZN(n220) );
  IOA21V8_8TH40 U36 ( .A1(wb_sel_o[1]), .A2(n37), .B(n79), .ZN(n221) );
  IOA21V8_8TH40 U37 ( .A1(wb_sel_o[2]), .A2(n37), .B(n79), .ZN(n222) );
  IOA21V8_8TH40 U38 ( .A1(wb_sel_o[3]), .A2(n37), .B(n79), .ZN(n223) );
  INOR2V4_8TH40 U39 ( .A1(wb_data_o[0]), .B1(n155), .ZN(n87) );
  INOR2V4_8TH40 U40 ( .A1(wb_data_o[1]), .B1(n155), .ZN(n88) );
  INOR2V4_8TH40 U41 ( .A1(wb_data_o[2]), .B1(n155), .ZN(n89) );
  INOR2V4_8TH40 U42 ( .A1(wb_data_o[3]), .B1(n155), .ZN(n90) );
  INOR2V4_8TH40 U43 ( .A1(wb_data_o[4]), .B1(n155), .ZN(n91) );
  INOR2V4_8TH40 U44 ( .A1(wb_data_o[5]), .B1(n155), .ZN(n92) );
  INOR2V4_8TH40 U45 ( .A1(wb_data_o[6]), .B1(n155), .ZN(n129) );
  INOR2V4_8TH40 U46 ( .A1(wb_data_o[7]), .B1(n155), .ZN(n130) );
  INOR2V4_8TH40 U47 ( .A1(wb_data_o[8]), .B1(n155), .ZN(n131) );
  INOR2V4_8TH40 U48 ( .A1(wb_data_o[9]), .B1(n155), .ZN(n132) );
  INOR2V4_8TH40 U49 ( .A1(wb_data_o[10]), .B1(n155), .ZN(n133) );
  INOR2V4_8TH40 U50 ( .A1(wb_data_o[11]), .B1(n155), .ZN(n134) );
  INOR2V4_8TH40 U51 ( .A1(wb_data_o[12]), .B1(n155), .ZN(n135) );
  INOR2V4_8TH40 U52 ( .A1(wb_data_o[13]), .B1(n155), .ZN(n136) );
  INOR2V4_8TH40 U53 ( .A1(wb_data_o[14]), .B1(n155), .ZN(n137) );
  INOR2V4_8TH40 U54 ( .A1(wb_data_o[15]), .B1(n155), .ZN(n138) );
  INOR2V4_8TH40 U55 ( .A1(wb_data_o[16]), .B1(n155), .ZN(n139) );
  INOR2V4_8TH40 U56 ( .A1(wb_data_o[17]), .B1(n155), .ZN(n140) );
  INOR2V4_8TH40 U57 ( .A1(wb_data_o[18]), .B1(n155), .ZN(n141) );
  INOR2V4_8TH40 U58 ( .A1(wb_data_o[19]), .B1(n155), .ZN(n142) );
  INOR2V4_8TH40 U59 ( .A1(wb_data_o[20]), .B1(n155), .ZN(n143) );
  INOR2V4_8TH40 U60 ( .A1(wb_data_o[21]), .B1(n155), .ZN(n144) );
  INOR2V4_8TH40 U61 ( .A1(wb_data_o[22]), .B1(n155), .ZN(n145) );
  INOR2V4_8TH40 U62 ( .A1(wb_data_o[23]), .B1(n155), .ZN(n146) );
  INOR2V4_8TH40 U63 ( .A1(wb_data_o[24]), .B1(n155), .ZN(n147) );
  INOR2V4_8TH40 U64 ( .A1(wb_data_o[25]), .B1(n155), .ZN(n148) );
  INOR2V4_8TH40 U65 ( .A1(wb_data_o[26]), .B1(n155), .ZN(n149) );
  INOR2V4_8TH40 U66 ( .A1(wb_data_o[27]), .B1(n155), .ZN(n150) );
  INOR2V4_8TH40 U67 ( .A1(wb_data_o[28]), .B1(n155), .ZN(n151) );
  INOR2V4_8TH40 U68 ( .A1(wb_data_o[29]), .B1(n155), .ZN(n152) );
  INOR2V4_8TH40 U69 ( .A1(wb_data_o[30]), .B1(n155), .ZN(n153) );
  INOR2V4_8TH40 U70 ( .A1(wb_data_o[31]), .B1(n155), .ZN(n154) );
  AO33V4_8TH40 U71 ( .A1(n1), .A2(n2), .A3(n35), .B1(flush_i_BAR), .B2(n156), 
        .B3(cpu_ce_i), .Z(stall_req) );
  NAND3V2_8TH40 U72 ( .A1(n80), .A2(n81), .A3(n82), .ZN(n155) );
  OAI31V2_8TH40 U73 ( .A1(n44), .A2(n45), .A3(n42), .B(n37), .ZN(n41) );
  INOR2V2_8TH40 U74 ( .A1(n85), .B1(rst), .ZN(n82) );
  NAND2V2_8TH40 U75 ( .A1(n39), .A2(n40), .ZN(n157) );
  INV2_8TH40 U76 ( .I(wb_we_o), .ZN(n36) );
  CLKNV1_8TH40 U77 ( .I(wb_ack_i), .ZN(n2) );
  NOR2V0P5_8TH40 U78 ( .A1(n155), .A2(n36), .ZN(n86) );
  MUX2NV0_8TH40 U79 ( .I0(wb_state[0]), .I1(n156), .S(n41), .ZN(n39) );
  OAI21V0_8TH40 U80 ( .A1(n42), .A2(n41), .B(n40), .ZN(n158) );
  OAI31V0_8TH40 U81 ( .A1(stall_ctrl[1]), .A2(stall_ctrl[4]), .A3(
        stall_ctrl[3]), .B(n43), .ZN(n40) );
  OR3V0_8TH40 U82 ( .A1(stall_ctrl[3]), .A2(stall_ctrl[4]), .A3(stall_ctrl[1]), 
        .Z(n44) );
  OAI22V0_8TH40 U83 ( .A1(n256), .A2(n155), .B1(n46), .B2(n47), .ZN(n159) );
  OAI22V0_8TH40 U84 ( .A1(n257), .A2(n155), .B1(n46), .B2(n48), .ZN(n160) );
  OAI22V0_8TH40 U85 ( .A1(n258), .A2(n155), .B1(n46), .B2(n49), .ZN(n161) );
  OAI22V0_8TH40 U86 ( .A1(n259), .A2(n155), .B1(n46), .B2(n50), .ZN(n191) );
  OAI22V0_8TH40 U87 ( .A1(n260), .A2(n155), .B1(n46), .B2(n51), .ZN(n192) );
  OAI22V0_8TH40 U88 ( .A1(n261), .A2(n155), .B1(n46), .B2(n52), .ZN(n193) );
  OAI22V0_8TH40 U89 ( .A1(n262), .A2(n155), .B1(n46), .B2(n53), .ZN(n194) );
  OAI22V0_8TH40 U90 ( .A1(n263), .A2(n155), .B1(n46), .B2(n54), .ZN(n195) );
  OAI22V0_8TH40 U91 ( .A1(n264), .A2(n155), .B1(n46), .B2(n55), .ZN(n196) );
  OAI22V0_8TH40 U92 ( .A1(n265), .A2(n155), .B1(n46), .B2(n56), .ZN(n197) );
  OAI22V0_8TH40 U93 ( .A1(n266), .A2(n155), .B1(n46), .B2(n57), .ZN(n198) );
  OAI22V0_8TH40 U94 ( .A1(n267), .A2(n155), .B1(n46), .B2(n58), .ZN(n199) );
  OAI22V0_8TH40 U95 ( .A1(n268), .A2(n155), .B1(n46), .B2(n59), .ZN(n200) );
  OAI22V0_8TH40 U96 ( .A1(n269), .A2(n155), .B1(n46), .B2(n60), .ZN(n201) );
  OAI22V0_8TH40 U97 ( .A1(n270), .A2(n155), .B1(n46), .B2(n61), .ZN(n202) );
  OAI22V0_8TH40 U98 ( .A1(n271), .A2(n155), .B1(n46), .B2(n62), .ZN(n203) );
  OAI22V0_8TH40 U99 ( .A1(n272), .A2(n155), .B1(n46), .B2(n63), .ZN(n204) );
  OAI22V0_8TH40 U100 ( .A1(n273), .A2(n155), .B1(n46), .B2(n64), .ZN(n205) );
  OAI22V0_8TH40 U101 ( .A1(n274), .A2(n155), .B1(n46), .B2(n65), .ZN(n206) );
  OAI22V0_8TH40 U102 ( .A1(n275), .A2(n155), .B1(n46), .B2(n66), .ZN(n207) );
  OAI22V0_8TH40 U103 ( .A1(n276), .A2(n155), .B1(n46), .B2(n67), .ZN(n208) );
  OAI22V0_8TH40 U104 ( .A1(n277), .A2(n155), .B1(n46), .B2(n68), .ZN(n209) );
  OAI22V0_8TH40 U105 ( .A1(n278), .A2(n155), .B1(n46), .B2(n69), .ZN(n210) );
  OAI22V0_8TH40 U106 ( .A1(n279), .A2(n155), .B1(n46), .B2(n70), .ZN(n211) );
  OAI22V0_8TH40 U107 ( .A1(n280), .A2(n155), .B1(n46), .B2(n71), .ZN(n212) );
  OAI22V0_8TH40 U108 ( .A1(n281), .A2(n155), .B1(n46), .B2(n72), .ZN(n213) );
  OAI22V0_8TH40 U109 ( .A1(n282), .A2(n155), .B1(n46), .B2(n73), .ZN(n214) );
  OAI22V0_8TH40 U110 ( .A1(n283), .A2(n155), .B1(n46), .B2(n74), .ZN(n215) );
  OAI22V0_8TH40 U111 ( .A1(n284), .A2(n155), .B1(n46), .B2(n75), .ZN(n216) );
  OAI22V0_8TH40 U112 ( .A1(n285), .A2(n155), .B1(n46), .B2(n76), .ZN(n217) );
  OAI22V0_8TH40 U113 ( .A1(n286), .A2(n155), .B1(n46), .B2(n77), .ZN(n218) );
  OAI22V0_8TH40 U114 ( .A1(n287), .A2(n155), .B1(n46), .B2(n78), .ZN(n219) );
  CLKNV1_8TH40 U115 ( .I(n43), .ZN(n46) );
  CLKNV1_8TH40 U116 ( .I(n79), .ZN(n38) );
  CLKNAND2V1_8TH40 U117 ( .A1(n156), .A2(n155), .ZN(n79) );
  NOR3V0P5_8TH40 U118 ( .A1(wb_state[0]), .A2(wb_state[1]), .A3(rst), .ZN(n156) );
  CLKNV1_8TH40 U119 ( .I(n155), .ZN(n37) );
  INAND2V0_8TH40 U120 ( .A1(flush_i_BAR), .B1(n1), .ZN(n80) );
  OAI22V0_8TH40 U121 ( .A1(n78), .A2(n83), .B1(n287), .B2(n84), .ZN(N419) );
  CLKNV1_8TH40 U122 ( .I(wb_data_i[31]), .ZN(n78) );
  OAI22V0_8TH40 U123 ( .A1(n77), .A2(n83), .B1(n286), .B2(n84), .ZN(N418) );
  CLKNV1_8TH40 U124 ( .I(wb_data_i[30]), .ZN(n77) );
  OAI22V0_8TH40 U125 ( .A1(n76), .A2(n83), .B1(n285), .B2(n84), .ZN(N417) );
  CLKNV1_8TH40 U126 ( .I(wb_data_i[29]), .ZN(n76) );
  OAI22V0_8TH40 U127 ( .A1(n75), .A2(n83), .B1(n284), .B2(n84), .ZN(N416) );
  CLKNV1_8TH40 U128 ( .I(wb_data_i[28]), .ZN(n75) );
  OAI22V0_8TH40 U129 ( .A1(n74), .A2(n83), .B1(n283), .B2(n84), .ZN(N415) );
  CLKNV1_8TH40 U130 ( .I(wb_data_i[27]), .ZN(n74) );
  OAI22V0_8TH40 U131 ( .A1(n73), .A2(n83), .B1(n282), .B2(n84), .ZN(N414) );
  CLKNV1_8TH40 U132 ( .I(wb_data_i[26]), .ZN(n73) );
  OAI22V0_8TH40 U133 ( .A1(n72), .A2(n83), .B1(n281), .B2(n84), .ZN(N413) );
  CLKNV1_8TH40 U134 ( .I(wb_data_i[25]), .ZN(n72) );
  OAI22V0_8TH40 U135 ( .A1(n71), .A2(n83), .B1(n280), .B2(n84), .ZN(N412) );
  CLKNV1_8TH40 U136 ( .I(wb_data_i[24]), .ZN(n71) );
  OAI22V0_8TH40 U137 ( .A1(n70), .A2(n83), .B1(n279), .B2(n84), .ZN(N411) );
  CLKNV1_8TH40 U138 ( .I(wb_data_i[23]), .ZN(n70) );
  OAI22V0_8TH40 U139 ( .A1(n69), .A2(n83), .B1(n278), .B2(n84), .ZN(N410) );
  CLKNV1_8TH40 U140 ( .I(wb_data_i[22]), .ZN(n69) );
  OAI22V0_8TH40 U141 ( .A1(n68), .A2(n83), .B1(n277), .B2(n84), .ZN(N409) );
  CLKNV1_8TH40 U142 ( .I(wb_data_i[21]), .ZN(n68) );
  OAI22V0_8TH40 U143 ( .A1(n67), .A2(n83), .B1(n276), .B2(n84), .ZN(N408) );
  CLKNV1_8TH40 U144 ( .I(wb_data_i[20]), .ZN(n67) );
  OAI22V0_8TH40 U145 ( .A1(n66), .A2(n83), .B1(n275), .B2(n84), .ZN(N407) );
  CLKNV1_8TH40 U146 ( .I(wb_data_i[19]), .ZN(n66) );
  OAI22V0_8TH40 U147 ( .A1(n65), .A2(n83), .B1(n274), .B2(n84), .ZN(N406) );
  CLKNV1_8TH40 U148 ( .I(wb_data_i[18]), .ZN(n65) );
  OAI22V0_8TH40 U149 ( .A1(n64), .A2(n83), .B1(n273), .B2(n84), .ZN(N405) );
  CLKNV1_8TH40 U150 ( .I(wb_data_i[17]), .ZN(n64) );
  OAI22V0_8TH40 U151 ( .A1(n63), .A2(n83), .B1(n272), .B2(n84), .ZN(N404) );
  CLKNV1_8TH40 U152 ( .I(wb_data_i[16]), .ZN(n63) );
  OAI22V0_8TH40 U153 ( .A1(n62), .A2(n83), .B1(n271), .B2(n84), .ZN(N403) );
  CLKNV1_8TH40 U154 ( .I(wb_data_i[15]), .ZN(n62) );
  OAI22V0_8TH40 U155 ( .A1(n61), .A2(n83), .B1(n270), .B2(n84), .ZN(N402) );
  CLKNV1_8TH40 U156 ( .I(wb_data_i[14]), .ZN(n61) );
  OAI22V0_8TH40 U157 ( .A1(n60), .A2(n83), .B1(n269), .B2(n84), .ZN(N401) );
  CLKNV1_8TH40 U158 ( .I(wb_data_i[13]), .ZN(n60) );
  OAI22V0_8TH40 U159 ( .A1(n59), .A2(n83), .B1(n268), .B2(n84), .ZN(N400) );
  CLKNV1_8TH40 U160 ( .I(wb_data_i[12]), .ZN(n59) );
  OAI22V0_8TH40 U161 ( .A1(n58), .A2(n83), .B1(n267), .B2(n84), .ZN(N399) );
  CLKNV1_8TH40 U162 ( .I(wb_data_i[11]), .ZN(n58) );
  OAI22V0_8TH40 U163 ( .A1(n57), .A2(n83), .B1(n266), .B2(n84), .ZN(N398) );
  CLKNV1_8TH40 U164 ( .I(wb_data_i[10]), .ZN(n57) );
  OAI22V0_8TH40 U165 ( .A1(n56), .A2(n83), .B1(n265), .B2(n84), .ZN(N397) );
  CLKNV1_8TH40 U166 ( .I(wb_data_i[9]), .ZN(n56) );
  OAI22V0_8TH40 U167 ( .A1(n55), .A2(n83), .B1(n264), .B2(n84), .ZN(N396) );
  CLKNV1_8TH40 U168 ( .I(wb_data_i[8]), .ZN(n55) );
  OAI22V0_8TH40 U169 ( .A1(n54), .A2(n83), .B1(n263), .B2(n84), .ZN(N395) );
  CLKNV1_8TH40 U170 ( .I(wb_data_i[7]), .ZN(n54) );
  OAI22V0_8TH40 U171 ( .A1(n53), .A2(n83), .B1(n262), .B2(n84), .ZN(N394) );
  CLKNV1_8TH40 U172 ( .I(wb_data_i[6]), .ZN(n53) );
  OAI22V0_8TH40 U173 ( .A1(n52), .A2(n83), .B1(n261), .B2(n84), .ZN(N393) );
  CLKNV1_8TH40 U174 ( .I(wb_data_i[5]), .ZN(n52) );
  OAI22V0_8TH40 U175 ( .A1(n51), .A2(n83), .B1(n260), .B2(n84), .ZN(N392) );
  CLKNV1_8TH40 U176 ( .I(wb_data_i[4]), .ZN(n51) );
  OAI22V0_8TH40 U177 ( .A1(n50), .A2(n83), .B1(n259), .B2(n84), .ZN(N391) );
  CLKNV1_8TH40 U178 ( .I(wb_data_i[3]), .ZN(n50) );
  OAI22V0_8TH40 U179 ( .A1(n49), .A2(n83), .B1(n258), .B2(n84), .ZN(N390) );
  CLKNV1_8TH40 U180 ( .I(wb_data_i[2]), .ZN(n49) );
  OAI22V0_8TH40 U181 ( .A1(n48), .A2(n83), .B1(n257), .B2(n84), .ZN(N389) );
  CLKNV1_8TH40 U182 ( .I(wb_data_i[1]), .ZN(n48) );
  OAI22V0_8TH40 U183 ( .A1(n47), .A2(n83), .B1(n256), .B2(n84), .ZN(N388) );
  NAND3V0P5_8TH40 U184 ( .A1(wb_state[0]), .A2(n35), .A3(wb_state[1]), .ZN(n84) );
  CLKNV1_8TH40 U185 ( .I(rst), .ZN(n35) );
  CLKNAND2V1_8TH40 U186 ( .A1(n43), .A2(n36), .ZN(n83) );
  NOR2V0P5_8TH40 U187 ( .A1(n81), .A2(rst), .ZN(n43) );
  CLKNAND2V1_8TH40 U188 ( .A1(wb_ack_i), .A2(n1), .ZN(n81) );
  NOR2V0P5_8TH40 U189 ( .A1(n45), .A2(wb_state[1]), .ZN(n1) );
  CLKNV1_8TH40 U190 ( .I(wb_data_i[0]), .ZN(n47) );
  CLKNAND2V1_8TH40 U191 ( .A1(n82), .A2(n45), .ZN(N387) );
  NAND4V0P5_8TH40 U192 ( .A1(flush_i_BAR), .A2(cpu_ce_i), .A3(n45), .A4(n42), 
        .ZN(n85) );
  CLKNV1_8TH40 U193 ( .I(wb_state[1]), .ZN(n42) );
  CLKNV1_8TH40 U194 ( .I(wb_state[0]), .ZN(n45) );
endmodule


module openmips_top ( clk, rst, int_vec, tim_int, ibus_data_i, ibus_ack_i, 
        ibus_addr_o, ibus_data_o, ibus_we_o, ibus_sel_o, ibus_stb_o, 
        ibus_cyc_o, dbus_data_i, dbus_ack_i, dbus_addr_o, dbus_data_o, 
        dbus_we_o, dbus_sel_o, dbus_stb_o, dbus_cyc_o );
  input [5:0] int_vec;
  input [31:0] ibus_data_i;
  output [31:0] ibus_addr_o;
  output [31:0] ibus_data_o;
  output [3:0] ibus_sel_o;
  input [31:0] dbus_data_i;
  output [31:0] dbus_addr_o;
  output [31:0] dbus_data_o;
  output [3:0] dbus_sel_o;
  input clk, rst, ibus_ack_i, dbus_ack_i;
  output tim_int, ibus_we_o, ibus_stb_o, ibus_cyc_o, dbus_we_o, dbus_stb_o,
         dbus_cyc_o;
  wire   id_pc_branchFlag, ctrl_x_flush, if_ibus_ce, id_gpr_gpr1Re,
         id_gpr_gpr2Re, id_idex_gprWe, id_ctrl_stallReq, idex_id_instDelayslot,
         id_idex_nxtidInstDelayslot, id_idex_InstDelayslot, memwb_wb_gprWe,
         idex_ex_gprWe, idex_ex_instDelayslot, ex_x_gprWe, ex_exmem_hiloWe,
         ex_ctrl_stallReq, div_ex_divDone, ex_div_signedDiv, ex_div_divStart,
         ex_exmem_cp0We, ex_exmem_instDelayslot, exmem_mem_gprWe,
         exmem_mem_hiloWe, exmem_mem_cp0We, exmem_mem_instDelayslot,
         mem_x_gprWe, mem_x_hiloWe, mem_dbus_we, mem_dbus_ce,
         llbit_mem_llbitValue, mem_memwb_llbitWe, mem_memwb_llbitValue,
         mem_x_cp0We, mem_cp0_instDelayslot, wb_x_hiloWe, memwb_llbit_llbitWe,
         memwb_llbit_llbitValue, wb_x_cp0We, if_ctrl_stallReq,
         mem_ctrl_stallReq, net70277, net70278, net70279, net70280, net70281,
         net70282, net70283, net70284, net70285, net70286, net70287, net70288,
         net70289, net70290, net70291, net70292, net70293, net70294, net70295,
         net70296, net70297, net70298, net70299, net70300, net70301, net70302,
         net70303, net70304, net70305, net70306, net70307, net70308, net70309,
         net70310, net70311, net70312, net70313, net70314, net70315, net70316,
         net70317, net70318, net70319, net70320, net70321, net70322, net70323,
         net70324, net70325, net70326, net70327, net70328, net70329, net70330,
         net70331, net70332, net70333, net70334, net70335, net70336, net70337,
         net70338, net70339, net70340, net70341, net70342, net70343, net70344,
         net70345, net70346, net70347, net70348, net70349, net70350, net70351,
         net70352, net70353, net70354, net70355, net70356, net70357, net70358,
         net70359, net70360, net70361, net70362, net70363, net70364, net70365,
         net70366, net70367, net70368, net70369, net70370, net70371, net70372,
         net70373, net70374, net70375, net70376, net70377, net70378, net70379,
         net70380, net70381, net70382, net70383, net70384, net70385, net70386,
         net70387, net70388, net70389, net70390, net70391, net70392, net70393,
         net70394, net70395, net70396, net70397, net70398, net70399, net70400,
         net70401, net70402, net70403, net70404, net70405, net70406, net70407,
         net70408, net70409, net70410, net70411, net70412, net70413, net70414,
         net70415, net70416, net70417, net70418, net70419, net70420, net70421,
         net70422, net70423, net70424, net70425, net70426, net70427, net70428,
         net70429, net70430, net70431, net70432, net70433, net70434, net70435,
         net70436, net70437, net70438, net70439, net70440, net70441, net70442,
         net70443, net70444, net70445, net70446, net70447, net70448, net70449,
         net70450, net70451, net70452, net70453, net70454, net70455, net70456,
         net70457, net70458, net70459, net70460, net70461, net70462, net70463,
         net70464, net70465, net70466, net70467, net70468, net70469, net70470,
         net70471, net70472, net70473, net70474, net70475, net70476, net70477,
         net70478, net70479, net70480, net70481, net70482, net70483, net70484,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347;
  wire   [31:0] id_pc_branchTargetAddr;
  wire   [31:0] ctrl_pc_newPc;
  wire   [31:0] if_ifid_pc;
  wire   [31:0] ibus_ifid_data;
  wire   [31:0] ifid_id_pc;
  wire   [31:0] ifid_id_inst;
  wire   [31:0] gpr_id_gpr1Data;
  wire   [31:0] gpr_id_gpr2Data;
  wire   [4:0] id_gpr_gpr1Addr;
  wire   [4:0] id_gpr_gpr2Addr;
  wire   [7:0] id_idex_instType;
  wire   [2:0] id_idex_instClass;
  wire   [31:0] id_idex_gpr1Data;
  wire   [31:0] id_idex_gpr2Data;
  wire   [4:0] id_idex_targetGpr;
  wire   [31:0] id_idex_linkAddr;
  wire   [15:0] id_idex_inst;
  wire   [12:8] id_idex_exceptType;
  wire   [31:0] id_idex_instAddr;
  wire   [4:0] memwb_wb_targetGpr;
  wire   [31:0] memwb_wb_exeResult;
  wire   [7:0] idex_ex_instType;
  wire   [2:0] idex_ex_instClass;
  wire   [31:0] idex_ex_gpr1Data;
  wire   [31:0] idex_ex_gpr2Data;
  wire   [4:0] idex_ex_targetGpr;
  wire   [31:0] idex_ex_linkAddr;
  wire   [15:0] idex_ex_inst;
  wire   [12:8] idex_ex_exceptType;
  wire   [31:0] idex_ex_instAddr;
  wire   [4:0] ex_x_targetGpr;
  wire   [31:0] ex_x_exeResult;
  wire   [31:0] hilo_ex_hi;
  wire   [31:0] hilo_ex_lo;
  wire   [31:0] ex_exmem_hi;
  wire   [31:0] ex_exmem_lo;
  wire   [63:0] exmem_ex_hiloTmp;
  wire   [1:0] exmem_ex_cyclCnt;
  wire   [63:0] ex_exmem_hiloTmp;
  wire   [1:0] ex_exmem_cyclCnt;
  wire   [63:0] div_ex_divRes;
  wire   [31:0] ex_div_divOpdata1;
  wire   [31:0] ex_div_divOpdata2;
  wire   [7:0] ex_x_instType;
  wire   [31:0] ex_exmem_dmemAddr;
  wire   [31:0] ex_exmem_lsDataTmp;
  wire   [31:0] cp0_ex_cp0Rdata;
  wire   [4:0] ex_cp0_cp0Raddr;
  wire   [4:0] ex_exmem_cp0Waddr;
  wire   [31:0] ex_exmem_cp0Wdata;
  wire   [12:8] ex_exmem_exceptType;
  wire   [31:0] ex_exmem_instAddr;
  wire   [4:0] exmem_mem_targetGpr;
  wire   [31:0] exmem_mem_exeResult;
  wire   [31:0] exmem_mem_hi;
  wire   [31:0] exmem_mem_lo;
  wire   [7:0] exmem_mem_instType;
  wire   [31:0] exmem_mem_dmemAddr;
  wire   [31:0] exmem_mem_lsDataTmp;
  wire   [4:0] exmem_mem_cp0Waddr;
  wire   [31:0] exmem_mem_cp0Wdata;
  wire   [12:8] exmem_mem_exceptType;
  wire   [31:0] exmem_mem_instAddr;
  wire   [4:0] mem_x_targetGpr;
  wire   [31:0] mem_x_exeResult;
  wire   [31:0] mem_x_hi;
  wire   [31:0] mem_x_lo;
  wire   [31:0] dbus_mem_data;
  wire   [31:0] mem_dbus_addr;
  wire   [31:0] mem_dbus_data;
  wire   [3:0] mem_dbus_byteSel;
  wire   [4:0] mem_x_cp0Waddr;
  wire   [31:0] mem_x_cp0Wdata;
  wire   [15:0] cp0_mem_status;
  wire   [15:8] cp0_mem_cause;
  wire   [31:0] cp0_mem_epc;
  wire   [3:0] mem_x_exceptType;
  wire   [31:0] mem_ctrl_epc;
  wire   [31:0] mem_cp0_instAddr;
  wire   [31:0] wb_x_hi;
  wire   [31:0] wb_x_lo;
  wire   [4:0] wb_x_cp0Waddr;
  wire   [31:0] wb_x_cp0Wdata;
  wire   [4:0] ctrl_x_stallCtrl;

  pc_reg i_pc_reg ( .clk(clk), .rst(rst), .stall_ctrl({net70484, 
        ctrl_x_stallCtrl}), .branch_flag(id_pc_branchFlag), 
        .branch_target_addr(id_pc_branchTargetAddr), .pc_new(ctrl_pc_newPc), 
        .pc(if_ifid_pc), .inst_mem_en(if_ibus_ce), .flush_BAR(ctrl_x_flush) );
  pipe_reg_ifid i_pipe_reg_ifid ( .clk(clk), .rst(rst), .stall_ctrl({net70483, 
        ctrl_x_stallCtrl}), .if_pc(if_ifid_pc), .if_inst(ibus_ifid_data), 
        .id_pc(ifid_id_pc), .id_inst(ifid_id_inst), .flush_BAR(ctrl_x_flush)
         );
  inst_decode i_inst_decode ( .rst(rst), .pc_i(ifid_id_pc), .inst_i(
        ifid_id_inst), .gpr1_data_i(gpr_id_gpr1Data), .gpr2_data_i(
        gpr_id_gpr2Data), .df_exid_gpr_we(ex_x_gprWe), .df_exid_target_gpr(
        ex_x_targetGpr), .df_exid_exe_result(ex_x_exeResult), 
        .df_memid_gpr_we(mem_x_gprWe), .df_memid_target_gpr(mem_x_targetGpr), 
        .df_memid_exe_result(mem_x_exeResult), .curid_inst_delayslot_i(
        idex_id_instDelayslot), .ex_inst_type(ex_x_instType), .gpr1_re(
        id_gpr_gpr1Re), .gpr2_re(id_gpr_gpr2Re), .gpr1_addr(id_gpr_gpr1Addr), 
        .gpr2_addr(id_gpr_gpr2Addr), .inst_type(id_idex_instType), 
        .inst_class(id_idex_instClass), .gpr1_data_o(id_idex_gpr1Data), 
        .gpr2_data_o(id_idex_gpr2Data), .target_gpr(id_idex_targetGpr), 
        .gpr_we(id_idex_gprWe), .stall_req(id_ctrl_stallReq), .branch_flag(
        id_pc_branchFlag), .branch_target_addr(id_pc_branchTargetAddr), 
        .link_addr(id_idex_linkAddr), .nxtid_inst_delayslot_o(
        id_idex_nxtidInstDelayslot), .curid_inst_delayslot_o(
        id_idex_InstDelayslot), .inst_o({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, id_idex_inst}), .except_type({
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, id_idex_exceptType[12], 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        id_idex_exceptType[9:8], SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45}), .cur_inst_addr(id_idex_instAddr) );
  gpr i_gpr ( .clk(clk), .rst(rst), .we(memwb_wb_gprWe), .waddr(
        memwb_wb_targetGpr), .wdata(memwb_wb_exeResult), .re1(id_gpr_gpr1Re), 
        .raddr1(id_gpr_gpr1Addr), .rdata1(gpr_id_gpr1Data), .re2(id_gpr_gpr2Re), .raddr2(id_gpr_gpr2Addr), .rdata2(gpr_id_gpr2Data) );
  pipe_reg_idex i_pipe_reg_idex ( .clk(clk), .rst(rst), .stall_ctrl({net70437, 
        ctrl_x_stallCtrl}), .id_inst_type(id_idex_instType), .id_inst_class(
        id_idex_instClass), .id_gpr1_data(id_idex_gpr1Data), .id_gpr2_data(
        id_idex_gpr2Data), .id_target_gpr(id_idex_targetGpr), .id_gpr_we(
        id_idex_gprWe), .id_link_addr(id_idex_linkAddr), .id_inst_delayslot(
        id_idex_InstDelayslot), .nxtid_inst_delayslot(
        id_idex_nxtidInstDelayslot), .id_inst({net70438, net70439, net70440, 
        net70441, net70442, net70443, net70444, net70445, net70446, net70447, 
        net70448, net70449, net70450, net70451, net70452, net70453, 
        id_idex_inst}), .id_except_type({net70454, net70455, net70456, 
        net70457, net70458, net70459, net70460, net70461, net70462, net70463, 
        net70464, net70465, net70466, net70467, net70468, net70469, net70470, 
        net70471, net70472, id_idex_exceptType[12], net70473, net70474, 
        id_idex_exceptType[9:8], net70475, net70476, net70477, net70478, 
        net70479, net70480, net70481, net70482}), .id_cur_inst_addr(
        id_idex_instAddr), .ex_inst_type(idex_ex_instType), .ex_inst_class(
        idex_ex_instClass), .ex_gpr1_data(idex_ex_gpr1Data), .ex_gpr2_data(
        idex_ex_gpr2Data), .ex_target_gpr(idex_ex_targetGpr), .ex_gpr_we(
        idex_ex_gprWe), .ex_link_addr(idex_ex_linkAddr), .ex_inst_delayslot(
        idex_ex_instDelayslot), .nxt_inst_delayslot(idex_id_instDelayslot), 
        .ex_inst({SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, idex_ex_inst}), 
        .ex_except_type({SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, idex_ex_exceptType[12], 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        idex_ex_exceptType[9:8], SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90}), .ex_cur_inst_addr(idex_ex_instAddr), 
        .flush_BAR(ctrl_x_flush) );
  inst_execute i_inst_execute ( .rst(rst), .inst_type(idex_ex_instType), 
        .inst_class(idex_ex_instClass), .gpr1_data(idex_ex_gpr1Data), 
        .gpr2_data(idex_ex_gpr2Data), .target_gpr(idex_ex_targetGpr), .gpr_we(
        idex_ex_gprWe), .hi_i(hilo_ex_hi), .lo_i(hilo_ex_lo), .df_wbex_hi(
        wb_x_hi), .df_wbex_lo(wb_x_lo), .df_wbex_hilo_we(wb_x_hiloWe), 
        .df_memex_hi(mem_x_hi), .df_memex_lo(mem_x_lo), .df_memex_hilo_we(
        mem_x_hiloWe), .hilo_tmp_i(exmem_ex_hiloTmp), .cycl_cnt_i(
        exmem_ex_cyclCnt), .cur_inst_delayslot_i(idex_ex_instDelayslot), 
        .link_addr(idex_ex_linkAddr), .div_res(div_ex_divRes), .div_done(
        div_ex_divDone), .inst_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, idex_ex_inst}), 
        .except_type_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        idex_ex_exceptType[12], 1'b0, 1'b0, idex_ex_exceptType[9:8], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cur_inst_addr_i(
        idex_ex_instAddr), .hi_o(ex_exmem_hi), .lo_o(ex_exmem_lo), .hilo_we(
        ex_exmem_hiloWe), .gpr_we_o(ex_x_gprWe), .target_gpr_o(ex_x_targetGpr), 
        .exe_result_o(ex_x_exeResult), .hilo_tmp_o(ex_exmem_hiloTmp), 
        .cycl_cnt_o(ex_exmem_cyclCnt), .stall_req(ex_ctrl_stallReq), 
        .signed_div(ex_div_signedDiv), .div_opdata1(ex_div_divOpdata1), 
        .div_opdata2(ex_div_divOpdata2), .div_start(ex_div_divStart), 
        .inst_type_o(ex_x_instType), .dmem_addr(ex_exmem_dmemAddr), 
        .ls_data_tmp(ex_exmem_lsDataTmp), .mem_cp0_we(mem_x_cp0We), 
        .mem_cp0_waddr(mem_x_cp0Waddr), .mem_cp0_wdata(mem_x_cp0Wdata), 
        .wb_cp0_we(wb_x_cp0We), .wb_cp0_waddr(wb_x_cp0Waddr), .wb_cp0_wdata(
        wb_x_cp0Wdata), .cp0_ex_rdata(cp0_ex_cp0Rdata), .ex_cp0_raddr(
        ex_cp0_cp0Raddr), .cp0_we(ex_exmem_cp0We), .cp0_waddr(
        ex_exmem_cp0Waddr), .cp0_wdata(ex_exmem_cp0Wdata), .except_type_o({
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, ex_exmem_exceptType, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117}), 
        .cur_inst_addr_o(ex_exmem_instAddr), .cur_inst_delayslot_o(
        ex_exmem_instDelayslot) );
  pipe_reg_exmem i_piep_reg_exmem ( .clk(clk), .rst(rst), .stall_ctrl({
        net70409, ctrl_x_stallCtrl}), .ex_gpr_we(ex_x_gprWe), .ex_target_gpr(
        ex_x_targetGpr), .ex_exe_result(ex_x_exeResult), .ex_hi(ex_exmem_hi), 
        .ex_lo(ex_exmem_lo), .ex_hilo_we(ex_exmem_hiloWe), .ex_hilo_tmp_i(
        ex_exmem_hiloTmp), .ex_cycl_cnt_i(ex_exmem_cyclCnt), .ex_inst_type(
        ex_x_instType), .ex_dmem_addr(ex_exmem_dmemAddr), .ex_ls_data_tmp(
        ex_exmem_lsDataTmp), .ex_cp0_we(ex_exmem_cp0We), .ex_cp0_waddr(
        ex_exmem_cp0Waddr), .ex_cp0_wdata(ex_exmem_cp0Wdata), .ex_except_type(
        {net70410, net70411, net70412, net70413, net70414, net70415, net70416, 
        net70417, net70418, net70419, net70420, net70421, net70422, net70423, 
        net70424, net70425, net70426, net70427, net70428, ex_exmem_exceptType, 
        net70429, net70430, net70431, net70432, net70433, net70434, net70435, 
        net70436}), .ex_cur_inst_addr(ex_exmem_instAddr), .ex_inst_delayslot(
        ex_exmem_instDelayslot), .ex_hilo_tmp_o(exmem_ex_hiloTmp), 
        .ex_cycl_cnt_o(exmem_ex_cyclCnt), .mem_gpr_we(exmem_mem_gprWe), 
        .mem_target_gpr(exmem_mem_targetGpr), .mem_exe_result(
        exmem_mem_exeResult), .mem_hi(exmem_mem_hi), .mem_lo(exmem_mem_lo), 
        .mem_hilo_we(exmem_mem_hiloWe), .mem_inst_type(exmem_mem_instType), 
        .mem_dmem_addr(exmem_mem_dmemAddr), .mem_ls_data_tmp(
        exmem_mem_lsDataTmp), .mem_cp0_we(exmem_mem_cp0We), .mem_cp0_waddr(
        exmem_mem_cp0Waddr), .mem_cp0_wdata(exmem_mem_cp0Wdata), 
        .mem_except_type({SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, exmem_mem_exceptType, 
        SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, 
        SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144}), 
        .mem_cur_inst_addr(exmem_mem_instAddr), .mem_inst_delayslot(
        exmem_mem_instDelayslot), .flush_BAR(ctrl_x_flush) );
  mem_access i_mem_access ( .rst(rst), .gpr_we(exmem_mem_gprWe), .target_gpr(
        exmem_mem_targetGpr), .exe_result(exmem_mem_exeResult), .hi(
        exmem_mem_hi), .lo(exmem_mem_lo), .hilo_we(exmem_mem_hiloWe), 
        .inst_type(exmem_mem_instType), .ls_data_tmp(exmem_mem_lsDataTmp), 
        .dmem_addr_i(exmem_mem_dmemAddr), .dmem_data_i(dbus_mem_data), 
        .llbit_i(llbit_mem_llbitValue), .wb_llbit_we(memwb_llbit_llbitWe), 
        .wb_llbit_value(memwb_llbit_llbitValue), .cp0_we_i(exmem_mem_cp0We), 
        .cp0_waddr_i(exmem_mem_cp0Waddr), .cp0_wdata_i(exmem_mem_cp0Wdata), 
        .except_type_i({net70336, net70337, net70338, net70339, net70340, 
        net70341, net70342, net70343, net70344, net70345, net70346, net70347, 
        net70348, net70349, net70350, net70351, net70352, net70353, net70354, 
        exmem_mem_exceptType, net70355, net70356, net70357, net70358, net70359, 
        net70360, net70361, net70362}), .in_delayslot_i(
        exmem_mem_instDelayslot), .cur_inst_addr_i(exmem_mem_instAddr), 
        .cp0_status_i({net70363, net70364, net70365, net70366, net70367, 
        net70368, net70369, net70370, net70371, net70372, net70373, net70374, 
        net70375, net70376, net70377, net70378, cp0_mem_status[15:8], net70379, 
        net70380, net70381, net70382, net70383, net70384, cp0_mem_status[1:0]}), .cp0_cause_i({net70385, net70386, net70387, net70388, net70389, net70390, 
        net70391, net70392, net70393, net70394, net70395, net70396, net70397, 
        net70398, net70399, net70400, cp0_mem_cause, net70401, net70402, 
        net70403, net70404, net70405, net70406, net70407, net70408}), 
        .cp0_epc_i(cp0_mem_epc), .wb_cp0_we(wb_x_cp0We), .wb_cp0_waddr(
        wb_x_cp0Waddr), .wb_cp0_wdata(wb_x_cp0Wdata), .dmem_addr_o(
        mem_dbus_addr), .dmem_data_o(mem_dbus_data), .dmem_byte_sel(
        mem_dbus_byteSel), .dmem_ce(mem_dbus_ce), .dmem_we(mem_dbus_we), 
        .gpr_we_o(mem_x_gprWe), .target_gpr_o(mem_x_targetGpr), .exe_result_o(
        mem_x_exeResult), .hi_o(mem_x_hi), .lo_o(mem_x_lo), .hilo_we_o(
        mem_x_hiloWe), .mem_llbit_we(mem_memwb_llbitWe), .mem_llbit_value(
        mem_memwb_llbitValue), .cp0_we_o(mem_x_cp0We), .cp0_waddr_o(
        mem_x_cp0Waddr), .cp0_wdata_o(mem_x_cp0Wdata), .except_type_o({
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, mem_x_exceptType}), 
        .cp0_epc_o(mem_ctrl_epc), .cur_inst_addr_o(mem_cp0_instAddr), 
        .in_delayslot_o(mem_cp0_instDelayslot) );
  pipe_reg_memwb i_pipe_reg_memwb ( .clk(clk), .rst(rst), .stall_ctrl({
        net70335, ctrl_x_stallCtrl}), .mem_gpr_we(mem_x_gprWe), 
        .mem_target_gpr(mem_x_targetGpr), .mem_exe_result(mem_x_exeResult), 
        .mem_hi(mem_x_hi), .mem_lo(mem_x_lo), .mem_hilo_we(mem_x_hiloWe), 
        .mem_llbit_we(mem_memwb_llbitWe), .mem_llbit_value(
        mem_memwb_llbitValue), .mem_cp0_we(mem_x_cp0We), .mem_cp0_waddr(
        mem_x_cp0Waddr), .mem_cp0_wdata(mem_x_cp0Wdata), .wb_gpr_we(
        memwb_wb_gprWe), .wb_target_gpr(memwb_wb_targetGpr), .wb_exe_result(
        memwb_wb_exeResult), .wb_hi(wb_x_hi), .wb_lo(wb_x_lo), .wb_hilo_we(
        wb_x_hiloWe), .wb_llbit_we(memwb_llbit_llbitWe), .wb_llbit_value(
        memwb_llbit_llbitValue), .wb_cp0_we(wb_x_cp0We), .wb_cp0_waddr(
        wb_x_cp0Waddr), .wb_cp0_wdata(wb_x_cp0Wdata), .flush_BAR(ctrl_x_flush)
         );
  hilo_reg i_hilo_reg ( .clk(clk), .rst(rst), .we(wb_x_hiloWe), .hi_i(wb_x_hi), 
        .lo_i(wb_x_lo), .hi_o(hilo_ex_hi), .lo_o(hilo_ex_lo) );
  llbit_reg i_llbit_reg ( .clk(clk), .rst(rst), .we(memwb_llbit_llbitWe), 
        .llbit_i(memwb_llbit_llbitValue), .llbit_o(llbit_mem_llbitValue), 
        .flush_BAR(ctrl_x_flush) );
  pipe_ctrl i_pipe_ctrl ( .rst(rst), .stall_req_if(if_ctrl_stallReq), 
        .stall_req_id(id_ctrl_stallReq), .stall_req_ex(ex_ctrl_stallReq), 
        .stall_req_mem(mem_ctrl_stallReq), .cp0_epc(mem_ctrl_epc), 
        .except_type({net70307, net70308, net70309, net70310, net70311, 
        net70312, net70313, net70314, net70315, net70316, net70317, net70318, 
        net70319, net70320, net70321, net70322, net70323, net70324, net70325, 
        net70326, net70327, net70328, net70329, net70330, net70331, net70332, 
        net70333, net70334, mem_x_exceptType}), .pc_new(ctrl_pc_newPc), 
        .stall_ctrl({SYNOPSYS_UNCONNECTED_173, ctrl_x_stallCtrl}), .flush_BAR(
        ctrl_x_flush) );
  div i_div ( .clk(clk), .rst(rst), .signed_div(ex_div_signedDiv), 
        .div_opdata1(ex_div_divOpdata1), .div_opdata2(ex_div_divOpdata2), 
        .div_start(ex_div_divStart), .div_res(div_ex_divRes), .div_done(
        div_ex_divDone), .div_cancel_BAR(ctrl_x_flush) );
  coprocessor0 i_coprocessor0 ( .clk(clk), .rst(rst), .cp0_reg_we(wb_x_cp0We), 
        .cp0_reg_waddr(wb_x_cp0Waddr), .cp0_reg_raddr(ex_cp0_cp0Raddr), 
        .cp0_reg_wdata(wb_x_cp0Wdata), .int_i(int_vec), .except_type_i({
        net70279, net70280, net70281, net70282, net70283, net70284, net70285, 
        net70286, net70287, net70288, net70289, net70290, net70291, net70292, 
        net70293, net70294, net70295, net70296, net70297, net70298, net70299, 
        net70300, net70301, net70302, net70303, net70304, net70305, net70306, 
        mem_x_exceptType}), .cur_inst_addr_i(mem_cp0_instAddr), 
        .in_delayslot_i(mem_cp0_instDelayslot), .cp0_reg_rdata(cp0_ex_cp0Rdata), .count_reg({SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205}), .compare_reg({
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237}), .status_reg({
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        cp0_mem_status[15:8], SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256, 
        SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258, 
        SYNOPSYS_UNCONNECTED_259, cp0_mem_status[1:0]}), .cause_reg({
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, cp0_mem_cause, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283}), .epc_reg(
        cp0_mem_epc), .config_reg({SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, 
        SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_315}), .prid_reg({SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322, 
        SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, 
        SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326, 
        SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, 
        SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, 
        SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_347}), .timer_int_o(tim_int) );
  wb_interface_0 dbus_interface ( .clk(clk), .rst(rst), .stall_ctrl({net70278, 
        ctrl_x_stallCtrl}), .cpu_ce_i(mem_dbus_ce), .cpu_data_i(mem_dbus_data), 
        .cpu_addr_i(mem_dbus_addr), .cpu_we_i(mem_dbus_we), .cpu_sel_i(
        mem_dbus_byteSel), .cpu_data_o(dbus_mem_data), .wb_data_i(dbus_data_i), 
        .wb_ack_i(dbus_ack_i), .wb_addr_o(dbus_addr_o), .wb_data_o(dbus_data_o), .wb_we_o(dbus_we_o), .wb_sel_o(dbus_sel_o), .wb_stb_o(dbus_stb_o), 
        .wb_cyc_o(dbus_cyc_o), .stall_req(mem_ctrl_stallReq), .flush_i_BAR(
        ctrl_x_flush) );
  wb_interface_1 ibus_interface ( .clk(clk), .rst(rst), .stall_ctrl({net70277, 
        ctrl_x_stallCtrl}), .cpu_ce_i(if_ibus_ce), .cpu_data_i({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cpu_addr_i(if_ifid_pc), 
        .cpu_we_i(1'b0), .cpu_sel_i({1'b1, 1'b1, 1'b1, 1'b1}), .cpu_data_o(
        ibus_ifid_data), .wb_data_i(ibus_data_i), .wb_ack_i(ibus_ack_i), 
        .wb_addr_o(ibus_addr_o), .wb_data_o(ibus_data_o), .wb_we_o(ibus_we_o), 
        .wb_sel_o(ibus_sel_o), .wb_stb_o(ibus_stb_o), .wb_cyc_o(ibus_cyc_o), 
        .stall_req(if_ctrl_stallReq), .flush_i_BAR(ctrl_x_flush) );
endmodule

